PK   �I~X;H)  h�     cirkitFile.json�]�s㶒�W^i��
� }��GUo3����S*�3�瑼��Ivj��P�,� �rC�3��"��C����M����׫����֛�j9��r:�l��W{��L'���|�������'w���b�ף+�՗���-�sJ��j�,\U�B��)��x�J�k!L+������O�WW���W������9'STB�B�V�� �6�ՎWZ��G���T�x��VB9[�\ԅ��L�k��[��:�HAZY{��,�न��)ѵ������B��,DY���M赮��֒8��+��j��m�̦,l�u�JZ�F��3��E����4ô,-��	ղJ��eT�:�2#��M�e�P-����N4��JZ��ꢲ��K�2]*]	��0:��J�"� ���Y?�DY+JNZSH+<\mC�+HEJ�WJ+ERV��~�y�J�W�j%oDQ��*�L��O{�.2(�Ҕn u�֔r �j�)� ���㉺ M��ѥ�� m���iX!u�vH�Ɛ:�!u���(��ML#E7��H�r$t9�� �ˑ��i�7䄒����i��M�\Ɇ�ƔM]4ڶ�hZQ+x!�He�V�\���S����&j9e��ZNY@���D�~D��2���4ja�D��H��h3^c��aD�)
.]a��f�5�kA4�R&�x�5��\e�a&D�:�20�y��:s�n`T�t�e���aRjh� ZN�W@S�r
b��b�u��]��'�۲1�hjn
Q{�b�*���8�$'b���z��UO�z�bZx`�1�ebԁ�O�?���W�5���_H�/m������e������l\D�Ҷ%��E�zD�.*p)iC�
�E�d�M%\Lࢬa�Fp)w�����eo��<�<����͔R86;;Bf9Q��Sf�&�66e���,�΃b��,���æC1q���WS�W9�1y��A1σb��<�)��<��YC�0�kt�˂� ��{k���',h?��2T�v;]ն(.��F���a�!�3�0z=n	C#��=�F��{�[��`�x�����Ac��4�z�G���Ü��
4d9�#h�q�G�H���
�k)h�o\cB�u��y�ՠA��]����	�e�B���и�a�^BX���:lk鞶k��aṰ,\x."�����Eg�b�p)�.x��/̓_��4�i�<�y@L��A1ˤ���A1˃b��,�Y�<(fyP���A1�dJ�A1σb~��������\�/8���r���KY��48���r�G��(p��l��!�q.����ACX�\�!,<��=��F��CXx.g{a�r���\����s�#������\���z��}���s�;�5_4NN�.�n3|��k��|�n�zr�1{�.�| &Y�1c�f87'�t%�$���"���t�!�VT��[aLj��'o�-�2D>�)����^�V�#Mrڴ�*�ղH�\z��&B\�~��e��W��*?�uIY�j��ZZg�g�e�����Ff�`b���aV	&��hh=`b�����i�I�T�@�1^
���K"��u�N�+t�]��0_����j��4�v����:���/R6��A���X��N��1�L�rc�����냹H
�>�ӧg�k���ޗ]61G죗����O�u�X�/�7��-\�Q��S�-�Q��o�-ܷ�)x/n\�7p�Fx�B�k�� ����^��w�!��}W��w�! :���/x�!���W�g�	��O�S�q� 	w	hOe A�=u �B��>n������;^ �� �_�P7~T�7��?o���byH8�^�����A�h��sd� �>C�'���?�s���B���id"A�]b�g�ؕ�Ԃ�T`�q9d��G�����:�b�K-@1X@����C9�H�.Y�`%_�U�X3��Ƣ�aQ̰(��	P"�EE�5V �e�&��c��Ѧ�L>Lpn L=��`0g��iB9��z�%�~p�@�]�� ' w6hFA�[J�@S��4Ǡ�ل�N6�u�u �,8���لQ�C�u�� �,83��YL����Bs���&-�:�p����΂�`��3��a�Èl=�8T��Sz�Ml=����tv��b/�HX��L�C��Y(	(����}:ya�hB$��߄P�����)8脀� c�x�9Æ�lP?ݲ�z�>:�vꢜ4��@߽��5X�;�`�5X��Bj�P��<����	5x���+�!�s�����"N��W��ƃJ�]mX	�;*A��D[*A��K%_�L�@C��_O;�/�6`���z�\pw>c"�V�����Ꮍ�A�6�NOz����rh��<껯�������,.�fh���K�Z�����q��8�+W�,b|/�G�K_�U���`�2��Gc�+�����*,2�b�t���K��������/�/��2����C���6�pŋպ)��r�x�M^pC��m� �+��":,b�"6,R�"5,��"=,2�"3,*�E堈>O��Ӄ�C���4"?ߗ�a���a���ac��#}�����e���٦Z�uHhiW��fPd�TB(UHS�B0�
��OC���qF�\�-�?�'o�������α���t��o��n����{�a�zt���u����e�_���v�]/����,��;�N'؇���_��ᱷ\�F&������_����N�Z��q�p�ֿ-6�������=-֮��m}�h|�˧��ۧ�[�	pLv$��QI�=���b�X�q���LN� 3�0��sB'��Um�j)�Z�:F�ͨ�eChk�e��b���e��
�L'���ϐݵ?yz��ź~p�9�XPμL��O��!�~�rV�;*�"Yd���c�,��Z�H&.���J�N��Q�!'E쨨��"AI��`ɶ���%|��C�<Б�ݠG
b!�MF�,61C��$E�b!㉾�'2R��Yl�#d���E'>BA�,�#�SF�LA�8��y�"��_%�E��(a��"�0F8���S7�Xl�>5��on��i":�3淭Ȟq�2�63�	��~<��3>��x��{D�u���u�ڂ�M$%���}o�{H�z����RP��K=�Q��ىJ���l����<�%#r�:2_�D9�G�~��ڗ����12�渙�L�}��]����/?�����_�����̿�?�TR��2�*��j}�YQ*f�+Z����M��7�R�ώ5-������? ���iO�V|���0��=��U�|��WP�y�z��Jd1-a�J4E�ͤ�ɍ�I+�^-B�ә��0���ޢ���0د��̤I@��h8�g��E��KI���W�*�� x徣Yj��/Z�W�^�bNGJx˝�Lp�u�y]��N�K�%�*��T�¶�IkZ���o����z����`м���'�`�2�G�*�AZOe��pBU�YyL%;�>3��>YװT3%�{*��
gbf%��Y<qIcYC�+ꠓDklQI��FH�j�e5�!�+�R���X��]A_UQq}=en#���v������e����dWVһŪ�Scf�˗�>	�j֚Zp?Ɇi�c��`�
Y	�lK<�U�CD�%y�����"K�u���r��K���?`�FL��=BOEg\���C�1:c�SS�Ehu��;L7)B�ׁP�ϡ,�GZ=-�]ە��IQ�3)�ڳ{����3�-�����~��s03+�����Ϯۼ<ꄜ	��������Pm��5?�d}X�������������o���������G��'�{@��~X,n����븹e3�vb�c��_�*�g���{\-��v�������~^��~�v�z��}�=���C(�E��i���(DN#DZϸ,�Yr�I(�@tF�P}�~?��ay#��|7�] �U V�WP4N�Ӟ�y��e����d���v��� y�x���"�Gi��}�<+.T��0;.Tֽ0.Dts��b��z0B���`D���#Nx�<'�XF���Y^���O�G��
��@l)(;�Uj+�Ϊ�c����P�] ݥ�=k��o\���,�Ӡ��*��B���e�d���@:$4ڠ`�~Yb+�ccH��hC�*'8`{,{)38�[��a��G�
JSC����M%s�C���&�\:,8⁛�怑I�������a��	,�/38H��L�[�k�Ls�R�#�Ϭn5����n5��t�ut>Oc$ ���G~�)�d� agC��,S��pv�xW���4��!ٍ��u�n��@�����b��eC�[C(?��P�FP�@���.`w/�..�f���N�g ��lH�Y�L]�9q��ٹ�q�6��q�qT��,eA�M��m�v��{��������d�!�m�v/�{���n
�!ٍ�t�ѻ�.�M�C&����������q�tWG߄N�<��{��,��~�s�xHW%�\L� �̀&q��j[0&`ת� �e�D ��.D��U��AL�3s��P�*.�����b'G6�T^�R	����K�SPR��X���5�쾾̰��@:$����V�"'�3aT1�1ȡ�U�H��bF���\D��=�}b�JP%ް�p���%�� {��D��W�a���5l�`�(��:�JU�Av��T)����9�2�=���
����n�9��%�f���kzd�䚐�xx����ݺ��>l&wV�����]�w�|�?����u_6�O��PK   �ZzX���7)� 
� /   images/0da2d01e-ca13-4f8a-b549-f8454ec0f5dd.pngWwT��.�v�2+W��]Y��h��˙"�M�� G����b��ܸ��l8��PP�'h.L����s�{���}�y�{��<��֦��9�cǎ�f����ر���}tߞ������cg����]����ݾ��n��Q�|p�S�_���}��;���/v��(<۱c����m�gnEB�z)ST�AF7��jP*�g�^{��)�ȝ;{T�n��u�������iƣ�xM�Q��;��Z����E��>���l�US�{&��h����w�n���Ԩ�+6�l��E�iij�����g���9�0ۿ�٪�ư��Ե��aq��B�85���p�N�����9�#r!����o߃9�M9�&��rK��K��x�����@?TV�Æ�]u�nKM��5�p�涾�؀�g��b����&#�*w���T5/c��>���h�K��ѐ�n�b��,�+�c��hUM�
SE�ҧH�q�@e�%�4�.̢�xgUT�U��Tg��\q�Y5d�����ڙ#52X�Z�I�@M�|t��Zc�
�	�#Sǰ�:���� �i�K��g�oJS��X�"fT����0�4�)����Z#��}sG1�1��2Wo"�ʼ1��%�}�Ƕ�����e:�m Y$������ڝ����bA��l�S�?��5����������A�l��A�'���*�z�02�W�VlV��)��Em"\�d����v^�6\�q��Cժt�6�e8�7��g::F:;~ھӐ����z�hZ���0�Ӫ�|cp��15Mî����?
�K?O�j�-�(��6��DS��`~Ԛ��[ʇ��:�P�!�-B��-�.���uƐz�:pҒ(�R:2R���aǀC)rAZԍ;�����Cȿ�o:��!��Ы�G����"D�;dT��[:|SIA���7_B��d$�����ȭ@�]���"6�3�g�m}X��y�����u�:��<X�Q؈(�~���1��Y���dW�މ&��(��J8
5_J�.}3"Ԙ���@�x)Qd�����Xe�f#�����7�Kc�Ѕ�z��ھ��c����pw����]��\H2ϿB������F����F�)N�(�
٫���D��r+x3|���m��I�ۂm��v[�ǎ�5z)�&��t���o��/Xx�w��]J<2�ъ_<�QyY~��v�"vU���)t���Vŧ_����hԗ]���*&=<5?*~� fk򉀵ܹ�
g~k���5�ֶ���򍲌W�J|��QQyUyJ����)5�Rո�8D�~+�,�}�X�(EY��ͱ�e��ѷ��V�����~�����|B�|Pޣ Hi���R�y[yG��9è�g����0��i*��j�f{�՚j�g�t}�w.*���4b�[��@�{�{��
����t>��]�H�f�V3ٻ˩�}bz����M=�J�m����|�&�Ť�Ac���зa<-4�n�;=�F>�ՙ{*px��["��Td��He߽��� gYM?Pu8r�.��Pr0���zo�m�����\i۾p��}�=��U2&��#��8Zz�`J�����-��B��������9��*������k����9��c�Q�^��?�9�F]��t��
����@9U&�*���ָ�C9�7-,�̚M�/}=
@z�r��w-Kׇ7��-$ M���Kx
v"d��I�/�%�T�v���jV��8����{��a��*P��%���鐩U3mY�Gn�g������� ��|��c�w�������ᶣ
����WX�RXl�O!7����8��s61.���S��U���kh�P�W�j�G�?��(<�a�U���4���#��|�����?J
�?��V2׸�����{�'_dH(������dm\~�W����SU�0@Y�]a� �/����y����ׇ|��l�la��F�++�8/��M��}U� @�3�z�Z&t�[[-w�4qP뇹�zo��#�A��6R��뷎����q%Q7N0�,-`��ɇ΂}����QwC]��m�i��=~��8�WY�΢���*��\�	�-���O�l�#�5�y:����m�;52����3�\��mRgq'��Q'���,���nW/)N]rpLg>~��*U6��*�M�����<`�R�������������s�{=�R��n]������Xj3�	�F����ڳ3�wf8��RN���7����׸.f����vs
<�i��|yL�ת�-��FexE���p&5��	��K���N��\�L%�WB"3�Z���)�_s�j�A�H�����0��4�[tv1;��1���
V�osQg_�n<�W0�O���Cݶy��.)_�]�.�:��0v��2�T؋���Fă6rj��W ~�o
��$���=d�1{�/a�m%U�P���8��\���]咽�*']��<�,���&�@^8P�b�,���n?�����\�/h��4HE`e���GS�[F������Sފ@xd|l��-=��׾�ѣ RP�����]�����F{ۭ����ak�J�3�m@嵽����L��%T���8��I%N��/��
"�fp���� ��z@yΪ��@P�KP��|���h��BgBF��~+~��Y��9��3޶�ŻCr˩�O�v�Al���eX'�4�\d�R�X��l�H�,��'
��}�O�g�	~ZEͯI�x:n��w��;`J�����]|N��sNafK���य़�����j.M7yw��DK����q�l�q������W%����οsZ��3�����ff�e�}ʺ�!��>�^�Z&�+��	L��q�ɼt=���ab�V��JB�TJ9���˥�u1�7� :��έ$�^ȱDV����H��u�}߆�.�_,`�.O #�K<.<*����Ww*v���3J�jj��F6�ꢲ��ҕ��!����b��%�X��.���#��]6���6�QG���Em��|[w[yAy��xnO�r"�͠]j߭G��>ٝ*6(����av�֣���[(�ϥ2f��>h^/lD�m)������9��k�\mЃ�m;~}T���] y;EФj�0�ǭ�?*YO+XQi8j	�?���:\*}��&A8����F�l�|���욹B~��9��R}�PIv ?Gs��!�,�
��;���F�x"4�8�z��k���+Li��%TQU�9�]*{W��1����
-�fw�&��ێj��+ʣ�c*��1���s��J�yGyK��/G>�H�Qe�Y�p^�E�pQ������4��d�1��+�{Z9�X܋���j�*񘜪�*�/�~�T��L���i��K�J���X)N�#O�Ni�3!���i�ّ����� \8Y1_b�$پs�џ���5�x���c7&-�B:5��y�g�+�IPs�	@���W	F�r�i�r���&<ۼ�6c�79����9W�|�>�da���^��NL�EG�����M�1��{�����;��_L��_yl��5���J����p�����q�� *��6�9̸:"�i���R��>_���]d�$�ܭyv}6v���:�C	�;�\a��P������P��������r�����g��%�p����i���b��ޥW�ׅ�U�>��pUxm�Q-�2�ƯY���`o]o��S��&~�C�d֏&-�B8-��|s�Y��qA�	[�,P�X��˧@�<u��٧���ܠ�m��l���6�t��~'�Gȡr��ҷ����N��S�4��}�K
: ���`�eD1��`�Z��:P�(*�bevo�b�I5��E0�heH]tK�w�]��HØ#qU$���3��[����9¶��q�1���RE�]ʠ����Լ]��Ƞ���1_x�0�h	����)i�h��%���/�ϡ�/��tGB��O{7�X������T��Z��8�����K����1B�l�#�cZ�5��'�e����c�Q�7��F?��[�n(��:�g���D��*|%Kŋ����;p��!xR��$Exk�`<a:@ݿ0�P��w�7���N$�5�*@TD>�u"���zS��Y�_���J��@����Q�{fE�N��_�9%�A�I���z%��� 24����U�Mm{t�J���km{ȕ��杭�F�n�R5���Qsqo���T�*�3�`HC#�,�	�q��>t���6A�+ٶ���Fz���G�I�� =����F�/�KW]���ƺxびJ�.s������[gI�Zdbad6țL��?��Ǣ��r��-�*��i@{��2'h~��[�b�i~�Vy�ƴl�k��ﯵ}Go�/�̽2�,�C��$�C�oOy�K���U�����C�����* �/��bҨ0R�x��bӴ677:�
b��	�(���7�kgv�V��n(�sW�|�ᓵ/c���(���Kx����u
1O�c&�1��FK�K����ϻ�ȶVm�᳂����#_! �J�[��0%��F�?R)��f���l��������>��W�ΩKAu��{��, �%`8����}�/���v8+��4��)ro�Q�G�se�T>���3�X*���l��t/O6
�1]uG{H}~z*��l�K��l���<��#��k����I�����g#��`�[��J�����T��=)�����n`�"��R�k�����yAJ��-8y���IQM=�h���&b�b��ǞbW}i�7�w��7Tk�/���p���2Z��۽F�R��$��5���D�R?R3��[~
��vd*�kr�T$�租Vݻr�ĭ@c��� |��r�-0���;�g��}��V.�����*P���5%���6'��{�R���v3/v�F)?��òB����������4��@lӆSܯl8ȫ��e�s5�[	��w�!g��u$W���;��v�`���G���DwQ�(r���³����r5��A��D:l2d�=���]��p�ӶOLӲ��.�����ڱ�D��|8��`�����v�:�����R韮ت`�h�Qd�r����0�r��κ�:�j�O����E��͘9����9�_�
��]"��uh���M)=�d��x��<�V�q��9�y�����r�r���N�gKs�G�?�-4�R�&2s��(��Q���2,�
�A���v�]�k�c����{�+�F�� �i�ts}��K���*xt���a��1Ѣ5<`�c.�qL"�]5�~$��dM�pd9i��ynd�~��@WL�$Um�����=�X�o�@��v��=�B*���Xf�#��p�T���0��.��'�������12B3#ݙ��g���VT���Ϭ����������z���Eu����\�V�=~5�k�J�%�#��#��2Ër�!\3+9`�&rӓ�x��S�@�j��D���ۚ���p�{�qG���O03n��^yjl&�jw<EW�2�
���_�nND_y���x×�%�7=���l�[�-�^ԧ����^a6�|��~���II�8f����r��m��ŋ��E��+��|H߬�я)s�� ���d�So?��$̡��b�&X4޷�Xĵ�pD�^�dT�C0�e�3�⧻�9�;�A��%�L\��N��|�͸ip��R4(�ăۓ
Gcߟ@�?
|���~�$�{NV,�c��1��6Ɗ)��bVM˱b���*4'=�y���ƨ�ޡ.�xֵ���imojm�1��0�-�ZWYd�QM����^��k���n��NU��]�r��s���[5���+�b|�&��5�1(�[1p|3�L.(�W!��u�\5�s�<N�۬�����*.�kbp@�1|��>8*Je]�z��"�8nޜ�� qÇ���(���9AO.�y�	�ж�
�IYb��)rc)�J�����Uc�
[p�p���#|u6�xz������<t���5{��J��N��|_Ͷʿ���q�}A�P�@>��0�Tܸ`��͏���PU.,~��A�W�BTU�������Z��QK�O�h�ύH�8��|�0��
���S�C�:V�_�x��|p @uMIգe-S�2�9���7���xVf>mZ��X�p(K(��d�3܏4���蚉.�cm5�M�u-,���KJ�?�Nxض��͘�.y�_��"���^���NBL� ɷP��Е���"T��"?�"��@j�P�ֈ��!dIHx�R��y�K0>e�a� �(�M-*v�eR�r�U�`�ۇ���_Ϥ*��l���/c�������r����w�}o�	;��Q��Q\{oн�hqo	�W��7G�îH.��g�i�Դ���Dw����	5�n�M��uĠ�쟗���5�=���[����hm���2�R�Q)�������_��R��� �M$qfb�@0����������UN�H;x�,��� �gߟ�l���!xO���	?�	��;,R��N�L��#i��K)�F�|;F�uؕ�]��*���=�M��)�Ze�_>�tڍ�FS��Y���>�6��O��OY���K#��Q�vS��xz�mX��{�.�>--��ڧr�2�ta;����k�f��� ���ݮ��k:vPݑ׶A�i̶�9!����V��VX�lZ��Kb9��@�m
������Aefdo4�@)N`]�tտ��=r��U{Hbh�Z���pTMw�{y�k�b,}����(Y�[AJm#��yz�z��v��������H��e�b�/�*�[�V��ߛ]᪔�-z���LGG��*�|lC�mP�]�&>V�[�ҟ���S��X�!9.T���U\��AFG[�п�\���M'��u;rcu����Vy������g���u����:�"P����`���'�r-���qm#b���/X��9�'gı@���KhЁ���;��Tw�t�
ཉM�����7�����2b�jSA?=�	�΀BI5N5���'�.�D�X���)�@�E)����-^����/xt����{p])�JE��J�Ւ������p�va&*�sff?�����]��K��Tzf�%E���˜5r�Q��el�ޤ[4xD�M�~Ճ��<g������y�s����Eg���J�����2�!Y��p�zg}���,\pC��1��m�
�z,�b�I����f���-�b�c6ڠ9���!�Y��hO�[Ow�9Sя2F/�.��Ꮜd���~nS��������=�Q���e���c%syB�runj�QQI��C\�__��tU*4��iZ2�Z��ǟ���/@\<�P�s����"(�C8^�F���Ǵ�H��
����WF�f�bH�mCwAFK��sりR(r:�KNv����c�Vͼ�̍b��l���O/���8��g��K����@W�l�O�UI���b}ur"��Y�G@!��G�/߾|��;�#㏚+�]����qT"�JG'�Ή�'��r"������7��+�va3�?|,��}~#��C�}�2le�M'dd�xf�RQ�c���e�\х�o�����-�FM� z�:V��8�^t��8vZ�h�<��_�Rfs8�W �i�~f�k�Y~7�TMP���WӉ"�'���ko����N�P$J�:`!����|�A��t��bL�u|n	��+'#��PeְR�Q����n뺼X���u��^��T/lR�5� L�"y߰��f��������)Y�jC��1��ם_&�EFLg:��`w��J����2�4�����erR�7d�-m~��I�P6��vl��i�v��!�7ܘ�K����Һ�vz|dwf�!�krJ?����.`������Ѱ�W��< ;lLzY�[�'LNq�t��l�C��d\�����,} V:3��`��|�i��Ӛm#���P��ӫ�}���w��=[��R��{66^ov�p�@�BT!�bAw$bl��v�6�*j$��KW�7L�Vx1�&�m�#q��_+�� �d	���{J���`��0�b���r�u��y�a��IGU��̄���\��PU#�L�@9`k-����^^��n��"�`�i윣����"<}����`6�����P �@��"*�*rG=�A�P��K_^.�><��;�-�����r(�т����Ǐ1����2ܾ�AT��3S��������yz����\�r�����ͼT����_E�z��0����!���~��&�`A�����O��������l+�p�~Va��I	`�E1(
��¨됖��\ ��>��%���f`�q6��R�ڛwQ�2�Ct�� ���,�AB4���/���&" ���nUa�m:�ڽVw�z:Rk�4��?��oV����a�t�f�e��j������_��z����!�M�e�ƣ[(B�߅�^�d@:A�S��ˠE��������Mf��ՅՈ����W<��i�X�hS�0^���7��gS�v�s�;���'>fu��Nv����� g�Y�ȸ]~��|�LBP�-���m��*ĝ�n�������}�^�������,�!���?(e;�sR������U�s=���u��f?W�{ک�`3��h�k6�M��z���Z^J��f�n�ׄr~>$��\��?�*Y%��̖��L��t�gj`��w�Vz�����״C�^�=�0�KV�����T���'¯o���T�d'����6!|�&`�� ��v�iBZ{�m�Yz�`{$�y%��B'��KEl�e�N��}ka��_��yOK��|n:Ƅ5e��$��@܃�kKl����+�c�s��o6�w!?ϡ� ���Gmݨ�xQ�>�I�z�S��X�"����!��W�M���� ���3k3���"�ⰽ�<�ş��ҋ.���>�B3P�۟X�us9�I�28͒�9@�P@�F��ZIC���:�¡Z��Dm�"_��9 L�@F�A��Y�zX
Ɔ7vé��<��\G�G!X�/����y�a-��i�5��f�Ƕ�d�C��H�a�I�፻� ��1?ֳ(>��<���ф�w��i�.�J���4�C�
Nt�`�l\E	�n�	3�uHs�"+z�+ͮ�qޡn��S��N��;���-��}c0b�.�n�Z��) �b���X�1	���N��|X�����Ո�)�mRg�,�އ�2;#D�3���pM����<��$�g��ٷ�9\W�,�;��uF��(Bi�&�ð��9c5N͏�6�_��g���Z�"1��ҐHu���av�v��Z{#,��8���\}`I��6�i������/�����,͊j�t�[�xw��A�f���&��g�����2�BΫ.�u�-��[��dC��
��u��X^��j=�68\��.A��ݍ.����D��ͱ|܏�UBqF���{��moI�B>�o%����C�L�/UvF�gu��G��Y�C�|���v�py�@-��O9W67t��il�|�8-an���s��J�sF#t�0^�QXD�On>~6V�U ����QCP�i�Q
o�1����v��*�M��N�jz�6��[�bW71��b���ej�J3.5n�"f����,�V�$tKI�����Dϟ8m��{{w�˚J3?�6O�_� 4.�ݺ�H��K�M�4�f�hxy���`����V�n���s�K@A���f�<A��⃧ 1�)�Ϛ�>�O+�\l8��{��Ǽ �]�aO�m_�k0��)�9��5B1�V�4���"�1�=�*ad\��p	c�i"�%��.���t:m#����PD)U�w`��������śd=�}������%Qu�HP�>ɥ�!7v�����@�j��&�j��z�\��. �� >���с��3�3�A�����O�A#ե��cݍ�	��b�港{���b�\Խޠ�R֘	
�����]�v�)�n` 5��*��A�#0!�	lI�j$��4��Us\LD��$3��j?6�fD��N4���WUWM��k�IM�BL��1��m�>��:P�!o�%�K	0�EB�5`�����թO��L8dF���T��"�	@����!�٦n}��~=��u;ĉhHX��'p�F&϶�V�Gt7�"ʉ��m�
�GB�����0}{���_^�;:��b�;mo�}�Z�y�^M\�i7�f�!�N�����%,8��[M�4)Y��d:�B�&�y��~G ��t�Ƀ��A�?�4[���ϬP��Y(��i�2���`��)4�>cL��1��D�&k�a��(yƴ��07��B6�n��w��UBR9/Z��G���u��-"��������K@� ��6<��˸�*5��+�^����.ǔ�-D۲���G��UbL��� N,MC��	V��[�4&,�h8�/Ӡ�@Q#|���VQ��k�O�=1���^9h>q6�hb�ꝓB
s&LtoBp�S$l��Ichi �����
�J�]��x�2n��*�W3��M�#А�B����A6�M� <�[8�N���8F@�2�y%�B�P��M���T��N,�h?�g�!kx�*k|a?��m�°�Py"�G�lM(��FO �Q��B�Q7 A���� }*����s�$��RՈ/'VC����G���� {jߩC����hxmq�3-U�`,�4�Q�
.��]ui|��gK��V+wڄ�]��7�)<�C>-�|B��h�+���E3>v:�E����M�K=�� �C"�:�;U1��)��~��\7���}�����j
�^�צ�(���_G2>)��<��j,�l����e]�|7]κk�U���oI�:�S��IDj�wh�5M���+�U���A(�*��s�g�-s��1ūX������WЇ 3�;�Ŏ�.Q,����~�>9�}����{��l�I���9�/�Gq��A;��)(Pp��iqW�|R�u��8 � \�h�{p�d��Y۰�%� D�h��;$���"�}7�<>�g�X��*ь�Z� �%�����2<:L#���	cV��uH�r��?�<��
��:!�MS��a��K�^D�	�D�]{02/_$#��!p�O����$�q���-zCm�:��*X���8�Ú�	g��d���M�����_ �~l������AJ	{]`ئNK�����������j��X���Be�N�@�܊��GR�B��)��`�6�1o���>g�n^T*�='�����o,�iG}���m?_7�1\���	5���,�T�t5���ǊV[G*d'��(�oX^�!1�1��TP=O:;fS:���G��i��Ȍ�B��R?���p�&�mV�j�f�7w�`����I��<m|��ul,L3 _����=g�W�3�fld-�]�;��ΰ#Q��	랠~��# ��(�ԋ�j��׫����x�sA�*��p�L՚��[�Um�D:s� 8�Y���`3�}�U�Î�c]gfdC.aщ��'��W	�ڜ 0*�_�U��/�?0k��j�9R��٘A5��JT�m7�2]�,K�m��S&�	�P�|n� ��5�$G�j�~�ͱ��"���̽2#&cۇi��[^�`M��Ryː�@�cE��uH`��h�������[��PR�d0ܣ= ��n��K� k��!�F���s�v�m^�q�ɓ�EF�y>������H���ɑ4�z���H� �Ax.�B�H%�#2w/�����n�	���Y�=Cb��{��x�3��n�$^�� �Q����aAU�#�M�*j�@���Lji�:�� #� [�DRis���o�<�;�z��L��-�96R �c�G�V/�}RE8�1vr�8g�h���4�k�`Ba~�	B���w�kЅî����S�b�ntl�3�������/��#J���ɵ�׮�;dJZ��>Pk��#��;t�ko�9A�MG�����9O�� ���"�#Oeƶ�k�O�t ����t~�f�ڏ]"X�=���N�,]4����.Q��=+w<%�7���EXkl*�싍G��l�/���}L"���#��|Z��C���F��'JY���ܭk���l>u)�����'�Y��%��:���!O)���� ���m>T��$�����T����g֡@xD�o&w0��w�i�n�3������t�;��m9��n�������"BږB���'Ғr{��0�(�!��m����w��9��s�''j��1���8Z��O��U)�[���ᚑN.���[ۜ��^�Q�(2��n�{PODL3Mϐ��=����q�����Y�q�IE�p9��>�%-��{-�mz�Q4�kʡ��[���ù��e|�Kưk�������`�����+��;��(��u���)_^�
3$�����5u������h�f�+:��@a6
İ��ې~S���sK��Ô�E��<�b#?�si��,�_+�g�j��@��&�b텎�.��O��5g�=�K҂�sw�5�wf�ְ�d�;��0I?�9�d�*�3S9^��YvH�Nڛ��9'���X���za�=}z�o|����l4&K9�r����{����k큩'7�2��֊�g�� �Clur���s3��%U�l0�8xɒ��̨�%D#�@�c3�I�̇��Îl�@~3&��N���q�0�7\	P(����Kq����eo���G�E���m�\�CA��B��q�%q�\�[�I�Ǭ��(v�U��A�J�t�"o�@��;ؒ��%^���jm!�t5�f���À�\SnQ���]Q���r��+yO����m�⾧��q�OX��mV[a��3�f=>z��	w�c��*�h��<�9��l��]D���<{�,|��9"���Ք��=���	sx�s�A���I��fW%(������@<���th�{넑�Gj����:5�"?���$i[�x�6hP�0s
(���|�g�������5�����h�'��8h�G�۟�w?��f?��U~k���/�zU$䷹0���9C�z:s���x��9�2�y��+m�k��X�ݗ�s����l{*�]P����W��sV7-��J�C�z��t�bT��܄$���s��߸ ԉ4�K�b�����sO�(P�F� 4�k�j�;��p��Ah��aR�qSdt�h�v-�NMGq.�~h^���{�ܙ�P3y�H��#R�l����}�Oy��%��V8�Ϛ�tif���kF����z ��D�Ly씇��c����*����}�!�UW���1z���%�?u���_~�ϊ�ˑ.~Y��R#�jьq�vfF��EL��A�(G\���W�گ��n�e�ͤf�s�|�Ls�u_�	��JW{��Ҕ�����L�>����ù�k���@Ĺɶד�ٌ2���N�ums��[��J#RNToaS���|ɼ����fBf�2]�-k�rĤ�*�ݏ�uCl@�+!�Q6@�Pp�7JJؔm��g������fG6�KϮ� ,ov?�f^N��
a������ G�9�O.8�&M�g#ɑ�"-#�<���	e��Wv���uK�!j�Rڒw��ڊ�,=%X͉+I*�X�P��#J볫��F����!a��ZU�t�F�OX5�X`������r�#HF��:�`�\2�9�����Z���Jb��~�.�kЊ�0A�G�݃}0��ɪ��A�9�`1~~������!G~DLg��W-V5 ���3"�6`�Z0�k=�Jb���[��9=�%xYz�oeP�,�y2`��	�n�e�����6B������dt�uz��
�	�s%*��GN���C�$���\�6�}�����)'�7}������[^;�q%3f�gpoI�)V����c��\�N`�c����_�0�4u��S:8�aByo)ɉ�됦$x��T\j�f34��qYc&J�x�_[֌ލyS^~tY�2`挸	"�P�@8��$�� '!� �z�����5 �4>��1Jn�Ci5����vp�с��z���O ��"S�<��D[h;,�_]6uX��\]��Ū�l�'؏8����HP	��B�l@�U����'����*_/8�NPnj����'�-Qk0wW�\��!���Iސ����m0y���b��?C�E>j�m(@.D�"|I���� Re���Z��Q~:bZt�L�O�X�������0�`���S��\�*���������ӠJ��}�����^���h7��{HU!�E~��x��u�����,�)��������e��F��s9K�����4{8mQi�.{dN�:X0K�% :m��,�g��� (@$*e��J��a������P�U�R��]5�*v�Nvܫ��Q����D6��Q�L�`o2����s>�;>��R�D��I�Pʌx!��U��8����;���k�*C
��]��Y�«��J���Y�;��!��X�&���t�kR��Om��˘��<���و�)���OJ��t_�C�`�lK�SG��{����Nz8���������*v֧A��rεV�� 9h��1�:��}��'�����̺۞Y������ ��+�b�t��#O�5�����\w�Z��[PǶ:)1���G2�� �`���v�"��r��k͇!%g����<��^�~��� �V8� �)&�!9�=ѷ�-��]��K�,���1��矮'~3$ �״[W��Z�YE�lr�z�l�7�.����[lw��N�2�f�A�pOp~�{�|��ك�t7�:��8gq5�Z7Dv��HN��5΃�[!�z�u����fb���k�t,2V,�K�4��j��RKb,y�<�}�$'	r%4��3Ձ=c��?z匹�,��z�bLkl��$�!�jw8�3G��G�5f4h�v�*���U� >h�NJ����I�>b��ƿ� #���;�I��e��RVXΊ��M�����z1ȃ���䏃��5S�������y��z��3���E�$���ү��/�D��o�M>��S��n\�w�*��>-�[1��D=à<����P�J�Xt���Zˬ�[_D��=ki3Oc�^������A�z���ҧ��p���W���V"o~>���l�Y�]FĔHuM�����9��1�vO����P�(˕Ň�@�j���Mg|՘�p�࿒]�ؗ��ŐZ�	�����_$��;��&Wp�ƭ<8�lR{3,&p~X�d�D[�B�Gc�͏s
K��N�o	����М��]n{ے��T����2�ᣬG;������	��B�N|�X��2YN�>%3<$8�rw	J��A+(�*f�E�UB�9 ֏i��H=��2��s;o�E���6��_�""c�?	�n�O�x&c��HF���:e��bs�ͫ�{eXd�1d�ύ@��K=n���1�㑉�x��{��(A����	��XN�&�u���P���B�,B�e���b��vp��p#
��� 
pU��tx�#�bM������4���-�.)�݉��Q��%�̢�Rx9z���[_��4���V���z��3K�L^繴:�?�a��U���r!p��e��zyf�5�#�7�/V�	F�&N4���Y��S����i�j苜Gu9�ܞ�NV����-�G<MT�T��xG��U��1��q�o�(?�3N]�Z]}��)�'��G��e��Z�ߓ/ɍP�+�*s����e�"�x��e�h8��i�ȿG5C��?h��z]u���5�Dv����X�Oy�i�g<��%$3O�7iyp�x�yݯb������tG���7��t'�ڶ�BTN�_0e�����Kі3i�ޔ��y�K�/Z���ص�R�X�S�efw_Sw�t{x�ў�Ꮃٛ�f!Gt�"�\t����L�lQ��"Y�����[Y��\"�N�&����v&}0mD/�$Gv���3-{�wݭ0���m�Ag�������k���;/[�:[\~���
H��f����Y�-�;n烝�N��zУ���c������������K!����QLyr�������������a�Ίݺ�%������;�;M���v�.���$������x�����҃��$��������Mw�����G��ٜpΞ))D�ew$+�:�����QG"e���I){����ߟ�����~�^�W��n@�/F%����R�~.az���d��o-�"G/��3��=�y��ȁ 8d����S��\JQ�vaƍH�un:���T?g��Mf���s�`��+����¾ h1�Y����bݸ��2�OĚ�.H�Mz���>��R��R{*EyQ����d�eBM0}sǭ��tx�l��S�I{�6kx�j>�Qf�T�(,�>!!�aNs7����u�n=��3AM��$������p6�~�(]'3����=��8��`	�V���6�R�Ї3X2@�Z��bx;)鄴
i�vL��]	��|^��g���(ks;�u��Чˎj�6Wqxo�
���Y�������}�����fYߣ"����������ozr�m�����z��/ʼ4e��g'�M{�aXE3��1�_?t�O��u�yn�ק*�w�k���ZE��;*��k*�۶�M�nQ���"�e��w���Z��$��}��1-���)��󏓫,�'o��\�,�<40�HbJ*�3��X=�@�H�S�i��"��`�G9����
���<�E�J����K^)g��g����xD�xpY�N�1ө��)�G�Wr;:v�Z�������;a;�
`�k.�u/k����-�p�b�ŧ��'Ȳ=G��3#�e��Ik�HY�ĩ��P��Jj m�j���_Ю�2��3����ؕ,
�zcrJJ��])�S�YsI�\�B[��Ʀ*���	 ao�S0,:T�}�7�z��%��?�t"`��o����g��O@WF�������]�$<q�۟1FK�谒z+@b�sR,�:��Š@x�
 R���1x賛9�ѩL�)���יOd���(cW�A�	�y�hGY���!w�lj�>�l 2D�k�zG��*�޹^�0������l�<p���y$�yX���CZ�(�^�tn},�J}l���W��%c��w�6T]�(����L�5q-y��a��ʖ;�����o�xh��$��OG���n��X8V��/IT�t��{�%ߐIY[n����h�^�����w`V��D2��y�m�����G��/�f��[0�gZ�>�V"��Z��8�M�˧i�^^�i}_=�y�V�䓷T���[�\ƃ����� \�?��K�v����oT%�qD�����i,R����#�y�V���{���&6�ds^�J{�|�
R��l����Ō_�+�7�$���t�Ń�X�)?� ��_fs>�LW�3�����E�z_P'�1c2@��w2'�E����@���eɄA+~��{��dr��ѹ��fz��0jh�fӕ���J��{Ys,V��	�Ҥ�i�������������<�AM�#Mw�(��ms7��Y�6Lx�G3l5��J}J�"T(�2|K�������Ͱ�Au&G/�!A�[���G�����ǥ��-���my^��G�*�<vR���8�ĥ�K�M?��E�a��z��U�gnW�x���p:`��z^]efZ����	��������'O,��˖l?���-g��\��y܊�K�� }vsԛ���W�IX/�j�ըp���Ir#�R�?���C��JY��ˬ|�2��-_\�_�O��M[�iI���jO��'��-����[Ѳ��w�nI^hu��k^+!�ʥ�K�-	�`=�Q͌k�D_S�WH��N���A��O&Yb��iA凐׺}q-f\~NM��+��(�u���S�?�?\n�ca��i&)RP��v�>Xw]F�J�|1�:bh���Κ^�ܓ�fǭ�b��賍yV�*�h��U��D�~�a��^�b7�ȁ�U�j��G0%��r�љd�1[�150z���ǲ�q?��EE7��t��cӚ�D��>P��i뎦㭷Ke��o��t���j)ۢ�uw�X�n`O��>MF^�x�)����Ϋ�287��u%�,|H�6�d���ߩ�����8n�#7���閮I*QB�j�����<�����	5�+-#�+J'c��}凪!?5�שׂJ�r�C���I]�})��I'yU���1�iH�6�]�ke�Ty�jB�I��3w�$.X��ߌ`��:jLR��(G����ǪY��L��A�� ��.���w�V�Ƭ��$ �k#��d1���}��j֝���dŲ<�������ݐ���}�w�z?�x	�]����b��$p�2sp�������=f�rJ�4<��~?��D�`���u
	F�]�Bܐ,R,	�2��[:y�k�z�������AM�����C����oo�Cs��&���J? ^�$���zU���'�nG�1�.	"�����H�(�4�ԝ�Ѓj�N�H�K�������e�3>��}����; Fw,��]O���nfe�N��-�y��$�	}��K$3����?��$�9��؜����|��iaӌ�[��&���-(���=��Kr4 Mm���~;��b�rk�y׎`�|�Iˆl�n$~.Y�����|���ּ��V�����[�$���*�1ވ[h�]�)����ѽ.�21G�{��ە��b��n���6�1���t�Na�'9���៰W��x�ح��7��g`P�w��k�"�����	�*]O�h�(�8y��!e���Z˭}EBK[�2��H��$$:����(�8�������ƺ*���+C^ 1���D�H�Lk��"���i���Ƭľ���e�jt��/�U���3��y�oy�E�ݎ�ڏ_!��yN�jv/i>��Wﲸ�U1 2$�V�M�m��  �ݐ��C�qP�����+q�[�j1�+d{�;5 ^}&�D_� 
� ]K�nl��dI<�7E�Uh_�3f���}&���s��|�g�Dʈ��p 4ٺu��`p�%��r����anL#�c�� h��@��Q��@	#mur�¾�I�)�cԐ�̨S��r�R`I����7	�l��\�&������I����v���0f)���6�Vy4+�Ķ�`��y�{D7�K,�����͡Z�*�� �c&FlS�m��C�Z�!zKMU��~у�*md�;�D�n!Ԁ:��l~��ǳWe�S���������b���G��pk2���2�'OԥLq`'�SĒ�ԕz\��9\]�ToR��hj�#�n���ҏ�;����e~��m��}3�3��Քvf���d�����,wRK&JGc=����e�t�j�+�aJ &��4�Dh�.�����8D��u���؊�;$-� ����aͽ�����0@~lK���#�|9���Ϸ�Sb8�"�ZR��O�E��1u�����A���c�OV]=қ�!�H�Z�A�|��/�A�[c�nl�ݽ`ߚG�9l[Qޜ���|��������zBs�E����f���^��u_a~���K��Ea|��Se<�6x�n��Б�m���l&�'#f��xz��ZZ_|	������<�������'�2s/��b��zM���?Ԏj�7&��h��W�ῲ!���l!7�l�d�mL�d�d�4��9����-x g�T����=�#���mF�-�M�}"J�f8�쨐�=�1\v�E�ZWw��0�����Ce�~Mk��/qg�황w�ĊݫD�Yp�cO�x�I�Q���V,Oq�R9f��P�%�4®e���5�)�|,+.u����)�>�;e���~�}�ռ���N�]�
����������f>�eQC'�b��y0w�U/j�bRP�3�5���J^g/�L��MzFw�����?˗ة4��a�ƨ��+�=���q/>G|��c����K� G�k�N�a�6v~���[�M�[�d�� ��,����Z��ь�n�w�Xv���mx$Ȱ�ƥ�U�%#`���]U�(u���"��v�����)��u�z=�+'�"�*=�0�;i&tCx���mP\��T����P�3�G�G�]�pe!p=X0z6T�RjX���Sr��z�i�&9\�lmpR|M��]��Z��X�HA�)�	a`�nƎ��<�n�ګ����*=�Q��M{�Kr1إ�*1@��1��w>��b��$q��{Jv�GI1�a��h�,bx&�}Ǟ�5���$��⮍.���D
�X���̿��
�]R��-c��V� gp�qM�����2ߠYl|.�M�#r�j��ϵM��o}
��ʑ��zQ��/��Tqz��,��"��M�?3��s�,!F�ű8�$������i߻����Zxi�S����f���夛�pc��^�s�ݻ�X�T�x0hﯸ�mī�)��6;���m�e?׆Q�
��k����
���6f/	10�Y�^�)(��n�]�I��7�`-�V:k/⵶ʒl?K���>ڸ礀^���Q�Z��'��NV/ӥ�m����."-�+o4��n�V�f�_m��~	>���㼴�Ң��7u⒧AH�����]�&���ӕR߾��Ï�m��؝����v�~�����܃�?�{�n'��D��u]Ú?T:7�m���t[��k�1������uba�{&^p�˧��0��T븙Tee-=����s��Hz��7T�i��GL7�e�M	�K8L�:�e����18�p��������V����(?c��
�|mJ�wѮ:FL"��_�;(�^A\���Ń߀Ȓo�G0�4�jX�S�hXԉXr�|%���0n�&K�Z�54�\����b�ŸA���WX4u��0���C���t����z����S�O�@�J+�IAEpG����+<�x1QS��F��02����'��
�
<�X{&�6��%�����u��l�U2C�������h�%��`~���S ��.�F3�Q�4Q�a��u`��HQq�=ԳZ;w���/����s���&�n?�L��ex�xZPj�--�臵Ɖ�b�
�-�V�8������SQzC'��Tjm��\�/b��F���x/ӄ�s��h�d�=�_�����"�q�a����"
{F7ןs����L(n:�T��E��d�����/N-x|/5&���V�7^����Yv���� 2�q�ua�Aq6��7R8�8"��-ݫ��/�)
�F�0�ԌFAK��u�?q���Z2�5.�`�#8E^���qM6T��F#,��i��"�gw��K�2'���r@�8�p�j���2�
�g�O!Y�,����C��&�x��^�[VK�JU���1�:�YR�!`��t$R�|'J'qGQ���u�~�R��d������p��U��`9��T{��x�@�/k���-8��k^�d����`���y-#�4�G/�=ݗ��]D&_��v�~|J±D�-���/g��y<M	��ε9�r��*Zv��\��D��:��{ΐ)x�kޮD������<lD�/V׃��0�&�v�g�9?;�تxz��;�:>��Y��Rg;o؛W��������<���S-��zt!�?�N�{o9iG&�;)l!�l�]�8����9ު���su(�{b����h���ڏ���ۮ#��i��=�,l��&5ߵx���Z��!T炴�.�VZ��I�$0�R�{�ͳ��(CrӴ��Il5�FP���Z�������s9t��dfB��g^�l�UeVfǢ3� �9�'�2j�X(5��&��5s4�mP�v9!�_>k�T%"�yB �DΨ���-���rpĠ{8y�2а�]cj0C���bkxq	�蘱��|�j$�o������,�%�����A3*,��YH�YI2�b�k�~h$��&7�LݎF�$�M{��-.��	PP���I�7L��0*����˛"��n� `�[p"�>�J���N�{�Y'W�x&�"k��9�,!�w�ʠi�KV�b�n��c�%��^Q�*�����ߕ�33t*!�z!�Ym�-^�����a�\,7&@EA��N�����c����d�i�@��r�}ܰi��y~�*H�󷡄�C,A��@�˸��/A�|�$*sk΍�C
we�c����fϫROmcKF[�>6�Tc�̩�ѽk��U[���ҸἜ^��^��u�+Og�Q�g	�cY�?����.�wEL��Rl�տ��|I��?3{OϹ�_�Y�!9�OV5�YЖ��[��\�,:[��%���x���({6$��� ��0V@�U�w/9��ZЛ�����U��p�\G����<�����d�HQ@����0_�����G%qd��BJbC��cP�|xG�2��$����z̙���,�,y���o�����5�˿��V���+��q7���s�y{��ٹ��ZO����@e�Ui���YM�q�Sڬ��uG=�QZ�����F᳘A�Na\CݻWl�1��f����B:�S�J�A��.�eի�7����/������'�5����(�z�Ҝ�P��xj�ב�()��4�S���H�o��K�����4N������r:3_��0���ή��D��M�<�<�f;^Xdڮ��K%��|�b���]��U���kz������*rw�mK�8�����d�%�l`<S&�k��/yUQd,# /+�Ջqi�����[4;' o�g��YX����:�)l��q,GYϞI
^��w�lm��`���3>lE��e=�z�4VT$!<�=����n�QE���A��ČI��9�����Д�8�����S�xo$B9�^8O��L��bO}X9k�,&�;�o��柗͵�-b��/ǁ��e?��Cv��^dJ�I8jz��,+��y*U��G`5v�t�?��=����6�e����'4̹f$�������+^[�C�q����Ts��/�o���&T0j�~gKJ9����߹��j���⢴���iN��'	o4�`X�-X�$����C�.�BlC�$�w�
!�V (}m�r�Z��s.��ۼ�?������"*���1�p���g��e
�w{�s����n�@wV��0�XU|�E#0g�lpc�"�/��Cf.�Y�mI7�q I��Eޞ�f�PD�h�eL�3
�8������z�}��뒹y�_Ъn:ю���V_�p����k�"��PU�&��]��]my�k?]�$����t���`{@��U
�l��2�*�UT�@�x5E�x�'�x�inb}Y"��U��X^q�e�c=Z(���@E�����j�cE��1:}}��P�8RD*���R�N�C]��$��ߢL�\�/׎��x�6�gҔ���si�u���I�aU��]o#�K��(��ƣ�R���_3�yo�X��u7�|G�ٙ��mڝP7?R�Be�䊲d�L�D벻u�˧�T��,b���J57S,F̄÷�������ZY��/Chq`���8,{�b̯���Ns(U�� ��� �bP����S�ڰ�%����/I��-�=}mg=qm�{��^j9`"�l_z�����ù�0�����Cw��y��|�^CzY��AEz]�`��=��)�^}$�����첄IB���7x�If'�߽��kR�Ԋ"���8Bc��x�	_���q�(m�5	����fN�B���$W��c&�x+������mڶ<N�RpZ#���0���I�AX.�����`t��ghP
����\w}�HN���s=;^�|�z�μS�|>�
��zZb��w�me���e�←FD0]C���S\�D`f��+��n9b��|�<Y�y��C��piY !�3��r^?�5���(2�1@�Z��Ӏw����5 ����$C����l�'����s��\�-ޕ���I������I�h�v�} /���K�]q*�\��?]��5&	�y�D͂���u��B��+H{0t�C�K'*�$D�� ��Д�I���l����I��n �I����8f�=ǉ;���#+����X3������%k�P�k�ne��Bڈ>t�x�Ӆ����ᵂ�04���eQ�gf�'��h���u�f�Է�A+�N�hb�[�g̰�"�!�\������M�.����8�%P���kਊ�2=\m����AmD��:������ǣ�U��,.�J��n5�>K���	-*RdD]}�pH���������p+�O��+j�ZG�.dg��s�X�PnN��*g7$������������{t��k������L� Ⱥ�B��.��O+$=�ڙ�g��J#�#n�tYn�C����4�:m�Y��BWٺ��
 |�[a���� K(�#�ƀ��o��r��x���XѶ�X�Ї�n��_�vx���C�t�Q�â�.��-�6 �ul��}�=�s��5���U�{�A݂�C~w���z���/6�3"�G8����6���/׿rj[������ۅ��|�-��N���z��4��B��SZ�^k)����i����К�ˋ���]Mtr\j�D��0U�u�CԤIKssJ�q�P�l��Nt��V�f���p�9��[�S߸�i��UuQ���3���dM랻Ԇ���k��ū\miE+	�h^�U�P���ge*�S�U_�]����U�\ЇjM��*}]F�;��o�殣ze2����gNc���	�����)l���k1%�x�B��3��=mZu����0���3{��t�����b��)EC;z�5���n�le�Ű��ŢZ �+�q>;��"y��0���i�_y}�Ȳ[���O *~{!T���.�K��q��҂g�d���nh:'�p�膡����1Ϭ��e�ؙ��Js�,i@6��,K��'õ*�q�7�Q,�:������������3�gr�$�(}[�\_w%�jh� K<�+�4O7��+qFt��sJ�P��LOJ�q����Ydڈ�V���&P��S���7�<eg
%���(N	x��Q�h����w��.��m"�(B4Î��
B*4��� �QoJ?C��*H��+�^�O`?ޏwc(,(k�}XF�k�������%�7����U\mȫB~�t��0�2+�ڃÐ4��������Y)��t�7r�z�[,H�^I�\�?�X����jU	}3@�y�芈XK��:���8�ԝ� 1@�=�7-~�It�.�f:C��{������|��!��s��m�t��a_f�D��Os�7ӾHy�L�Č�U���XH8Ct�Y���ܝT�p؜ ��(���	A+%��x=��1���n��s֐!�75|g�b��<��R���x)��J�2&O����{���������ҫ����FXH!^_G�ge�]r���=/I����u�쾙�(�O�%yZ[��N�מek�ٿ'�l�&�m'��E����x}��jh�W�:gK���dj)� �Bme�Ia���!�c��R��-��+o�1�� ,?�'��*�����a������?�Э/�,���ɲ��X%(xs j��R�eЕ���8�U��w8إ����	�E}�֬3���������(� ��ګu-�j0�T���� ���n�d�a|Іy���Q����^Uͨ�RV�u����G�����BJKH��pG7a��x6�!CF�
J�-x����>�@f�����M,�l�X����	�5H��z�<T�����S�s�`vҡoaד2Y�����w��!.���c��$=���5@�n�B[�����w���r�8 iDM��!Y�yiJ��F��Q{^}hF;p|~��2y�����ݫ|��ʼd�UT|5�&�h5��'�ٯ!��\6�*u��E�xf7�[+��V�P�{y/���A�B�
(W���7�� �����hU콖��H$@x7{U�L��^0:"�&�(PUD����2[�������P�oi�*	�M�/v����/y����P<s杬c�8��ү_�I���q�$|��X���Z���\�	A&�^��ۯ�%3���b����%-�a�^X��(��}WՀ^j+� �i���4W +��w��F+��6�Ć��6����-��̸8y��M։�vzh�u��uk��q���/�mu��y��}߽�|ߊ��e��q�c��S)�Ӓ���^���j6����������e�,iJV2�ٲ�~���x9���I�E�'ǿ}x�ŷG۰���^p���0ܙ9���v����-��o�w�k.�/��;���-����� @�{����|��~�2�7� `$�jRoo�O%R����ߌ;��5�N	@�f c�����^���+[kN Ú�;�?�[���3t����Z>@��x����j�j��/�L�Z�;�E}+)�$۠�.lV]ca�����|p8����?Gt�L6�4L��8L9�� i�{?E�|)8��� :\}�"� F<ĀҸ/�j����3!������4�7�,N0�j�s�%S�1z��؉7���r�YF_��u�2;ٟ�`�YH���?�sK�/p�Cw�]Ob���%�3W ݢ�Ht��T4�����C�w�5�t	�����$���-�Ek��Ǘ���ۓo���CEYM�n=��)�Kf/�§)�D7�����Nl�Λd'�ߓ�3}�	@U�#R�Z�!$�����LC-�d���X'R����Q+�*��+d����Ǭ������8 �W�RvǮ�&�h�<�Տבؠ���}��t6ЖAJ{ϭ~�3$E�Ip��{_#Ain�d��=�M�V�����׃%���&3wC�j
�����{��0�u��-G;Ec(�l��INS���t|�@i=��ق��;�_��z���A�C{[��|wM�LN���3{�}.��e��%в���o�ݕ�!'W�o�zkg��MN�ZӃ�f�$����?�<�=/�K�?~�>���ꏋ��'�����Yc���&S����hJ*g�����M�K�[	)L}����kS��� �P�k�6T�u�֚��u�9�Z>��	�jˉ���A�~�{җL�^Y��n�[��z��dV�������Wê�ܯ)�*61��/��2����F��c.��.42��y�O��0�T�R��<��+����d�pCOq��-jq��y�Y��4��$lM(Q��Qhoa���@l\���e�CB"���Oa�܍N�uĂ���F��J�p&z��N�w�D�vb��K R�"��w���6B��NM1�U vʚ��F�%�dc�]��؅�hq�!��M��`P�(ٗ��t��}U���Jw�u<F���H�G([�}�`��] �t�Z�R˅ ���EH���sy�8�Ue��3� �}9+�d��T�+�Y�ĹC\D�j6(}�d�1C�a����������j��k�Yz�L�-��q��x�(r�mnyႲ�%�*T6Ò���/�[4�S��5i��WM_�z�i&ހT<,�7�	���f_��T�HAr�@b�8`E��*Z�M$XW@A?���C��5t�u\�r7%[{�ՠ�@�� T�`.�ޘe��%�� J;�&�V:Zr}�
��ub)>���e k��}��Z1�lw�G]�{-B����0�2�V�DI
��v#�� �l����L=c��Oۜ��Kj��m�3 ���p}3ҽ[�{)O��������Y�yB|!��^`%=��U��gy�i*vCz}s"���kb��h�Y�V��G_����z���wg|:�YfV�ڷ���\s�������1�w�BO��ORC�7 s\��T4�y�ϩWv������͟���p���œ������.^�n^�����T幩y6}eh�0P��1V`������K,����z����{�Ɇ~˪��}QK�9J3�Zk
�������aϐ�^����O9�;e����$�~̷Ki���l���O�t����SkK�'�v�õJ΂k�\Rp�z`�꣣]�ad���wG(� ��ۍ�1G]��ӟ7M��$����[mf�ņ�8�hD�9�dW�Ě$�B�Uӭ*p�kȤ��#k��b��x�2���p��D���b �,�,BkTg�*�6���\����K��k�n8l e���4��AƜ��Igx#*�VR-� /�HP,��-���ؗ�+��<~'�z�������R �j2��.8��� t�'1��Y�R���*1ڢf�$wQ|���Уe�đ������ߥ%�vo��8���9��qvײ�J �E ��]����m�]�%���T;0C�*�����W&=��q7wJ[������M��٬G�tR�g�*��P�2�S����MW���g�;!���䖲�>�Y�����w7!$(� ƀ:������/�0���m�	�H�ڟ��VOZd����T4Z��qf�ȕW� ���ኰ갇_�(�Ho�0:�@Q�[ l�����������P�-�О��b�����!�j��6���*My�S���G���j�V�.+��l-�w�Q�Lכ��_��l����k~}���C6���%ߞ��̓�\����r�{5�<nU�cd���Ky���PUZ�v��
zLA�o�-L��>�H�Z&�鞻�	e�|�����t��7����
[��w^KU��6�Nq`��e�����	���ҡ�RE޾��*���a0Rx�]R	�Ϗb[4:�\2��<���?�t]�d�A�= ���3}�&�kS�U���݅/���@�+�s�Q8nH���bS*��Pi
<���!�F֐D�c|�4ع�A��0悏�r���	c!˧(vF����g&M��p^�A�ź���b�����a�!C������22����DV���o�����$��H���ш�8s@� 
`;W�ggzZZ"�^F\K�r`�&m"���m�p��X��
z��`�1�����+l쌀$Zrw��@�NH�ZR���[�v�AU!xo���LI�c9�6�U�*��E�~�w��� �	"&o�y��Xkvخ��4[�������pzA�D§A��ھ�ɗ�� �BlsC�W��C!����P��-�Ffߪ�lx
���wL�� /a���%���(�4��oU��4��g)h�Bb!����v�:J��x��Ao얣�$���?��/(� ���"�3��[o���*��K`�ڠ����]Ͼ�d��ʁ�8?L0x�eax�%L��J�~.\��Ff�ˌ�f�����s��D�Xy����nB���y�uӳ`�����Bp#=�>����r�T�� ����2��_Ae_�����wf�V��7�#o[I$��^z[�����n��Ɔs/����DyX�K؃�3U�'P�������`��Ë�agҏ6�w�O�^X���&�'���p���.I�P���,S�W\˭	L�C��?��/B�(� pD�A��A��������CM���O{+��k�-�~�}_ ��Y`��7GI�̷��b��h>B��M����&�[�Wm�ˢ`�S��؋�5�en!�cLV��[��(sZ�/�ڮj�%���.��@�U�آ����*PjU���g@H솯�r���*S���F�q 9��(�-l5�X"�	�aWٕ���p����4:5��a ��H���]�~���x)����K���,��S(���n��w�Pwн��p�N�F���h(��4�jp�)��Ĥ8 ��ǂ�4@��'07@��ȂjY�:4��X����"�����-�s9mb)���h������f�Qh ,,kY���0��o!�{�o�O�0�=P��=��Ŵ
�H�;x��>	������h#,rx�O��h��8e�������_z�o����T|�IG ��!����y�F�NooE��6���#�k�p3�@+���47�D�ǯ��$�d���բ"�����7�\2&�ɼJ2p7��}!tl�nբ��_,K�E'-q�u��ߺ���.�XZ)Í��c�e3դ���Kf̌�C�gy�������Lݻ=��D�&�Y߮�9���'��߼�f�b���u�ebk���z��������2�hۂ]m��-&mk<mac>No}La������OH�w��2��j��O�.W�ܲ
�����~pxV`�w� ��Pj������ʗ����䆶�]��*�$k���omiz$�*B�>�nv�ixM	1���/&�DT��8H�5�t�A����	"��&��"��Pj$�fؔ�aKs�ų��7�y�8P���Y�` �Iح�AMQ�Ĳ�r~�������d�z�=q�y Q�:i$Ҋb��~��b7�z��xt�)	-��#�o����!�S}{5�����r��Zn*ϣ��j����,��� �:�:>�w�x���&���N�9_�2�C'B�D֦H��$QQ캗N����'e�,L~�)��S��[�L�(�~(̚jgUF=�0���1�hf ��D��������bw[$L�������k����Q3��995���z��$��G�^Z�t�;{&轡�aӽ�]�ty@�%SK00;-��ʿ�[eHڲ���J�*�r7gmČ��-JH��뼲�e�X1�p ��'zU�d�e�BYk1��?)n(�1�wW<�ӰS�1����Kh���$"�"�z��?m#A���ri��?i�6�گ���r�O~�\¬��-��?����k�vw�g���_�U�$�SD��d�J������b&�]%�G�{��`��h�Ag����jqDS��#6�I�?$j��i��ZF6�f^cY��@�� 	��wA	ᄞ��sD7���J��,���.Y��>-�L`[[u=8�}{;�"Ѹq���U��;��N��ܿ�~�"؟�ē�ݾ���z�+ì��Y��d+��X��)��kIIv ��5?�ύ�y?�_���ɖfu���3I��$�_$M82<���կsfdܫ��������L��k٘���a�a��~�0
 B��C�A�zZ��v"5|@�r�f1b�0���M��U�it6�~ޏ��x�{C��V��#���S�F���4Y#g��l��y^���K��em}ڿ�!'�wU�c���F#����X2�D]��ĖEg}�WA���I�c�3sRa�Ɯ�]���Qƌ�r"����7���Þ)��r�, ⣓�Yqـ���� ��랴*�ا_&@�O��S��F�.z 8�@�tQ`jR7W�%2�+0ާ�1
��"�+Q^(l�7��O0A�q!�{[�����P7}��R��(]Z*޴c2�׆@ƈv(��
������"HL��C�ؠ�Ul�c b,�8�Xo4S-�3*N��j0��؁ʪ��Z���1�w�E�G?�Q`�Sq��1��o�K�R_�-CѧܙĎ��j@c���W0W�H.�B��1���*�c4�OB�Tm�tZ�H�%=�jɉ^�7���A��n���Y`m �諾�8,砖�+4��o�zw(6ɺ5���yJGJ�3	��&8�JBl����'�P.ʷ��\F>��"@��q�=�s�<���G�}�cUޓ��У���s�T7�,�gkt�-���P�t���փP��4)`}��V��D�K��ӽ��#H��q����}����sh�Ѓ��%�1}��:,#��ߛK�:[�仐���Vη��P�/˒ه8�2&Xe����Qz=|P�}�''��]�^�I��z�z\�b~���3��:&׾�ES�P��m�^��/����x��UU7B�NYԏ��喰���	V �䇵�<��m���y)��k ���2y�ܸ�U����T��Q������u��� ��Cx�E�QG1$S��AvF4ي-���Y6yU��,�)�p���gWB&�%�@�s��Bk���F�!O�*P����x�����(��h���4s�x��	�{I��!�P�"ǲ,�k����`~��F?B��T��r�qz��z�U׻���4�88���n�,i1�g]Iƙx��Qc!��-5��v�W|TG3&]r�)���ٽ��8�_���b:j��I/��>�I���:�:�v����i[3���"���N �����6wͯ�-��'�����6 �?��l^�h%�z�sz�?�*�"��$`��<����wy՗:8��by�v��5x�@_��5\w���Rj�T"�S��*��x�x������B����Ӹ���KR����p��Q�L��&`������C2T�]IT�6�JJ�1�F��z�ٹe��/n�դ����\����8~va3�m�s�\
��b���f��B�w5�K��HR�)�Bn��;���BnE��.?�?�<���y�^���s�"i�Jc��6vL���?�����!��q>A<�W%��w!�5澒�7m�[Н?�&�U����W�V�������q���y;�{�!L�(��P�)+���z/jk"�|Q�n.Y,N2�����<�����10Y����ټ�6K ��q��ԉ_��Q�05	�m7"/d�����Y�	�:�����[VH~sh}4d6Ԝ�tDz;¿],]j�;��t�6�f]�j~���n����
*��=��2oڈw�in~�1v�s�-r�2֒�4����-��-�ן�]�7���N�N��F/=*���K��M^7Vf��\���[=�����2��e������{��	������-��}�9�":p�!�nx|�f��\x�Zg�K��#��ϳ�b��c�M�
�V�x��� )8-BJ�+)���S��f�S��h�xfy���Ǝ#}�1n#��1��c��[���h"}��� l��l,FG�����X�d;Uoepjo�Ib�MD�]�֊|�G\�#��S5���E �>(� ��X���0�h��E���/�xKq�7E��ڗ;�7;����߃E��� 9��r��E�Sl�Y�y�@l�Y� �4� ����o��!������9�Bg����D3�	�8�N�Qh�L���{��b�4��>vfЧ��)ڴڮ5�`v�C9^p��^/��o�l�i%��]zHW��G׊�ٮWn��7f�ST>c(�>�����)�Zt�|\���>y�ٿ�1�ː�W�#�G^V"}����8y"[r��t�����1WF�"J�'���\J&�����W^j��Y|+JT��QX��YKAM���������Ԕ�m��}��)_��~������m��g)>��Y�tF�Ja���\��
b�qQ���E��,w��˩ah�X�͒��n�Y���p����C�N�b&mU�x��Rz@�k,�1��b�J�G�W�E�&N�H�G�<x��L+��5���0�����.|S'�N�JoxP�k=��&�}
�D`�(w<x>b�\"�Zge���R��j��_y��z�e���9�Oo��k\�ql�x25�?v�ݱ�N(~%��r�>67�ܘ+k��,{Z׋�}�a�ky��q$N�.����u���ڏ��5h���$�L�Sb�	�n�c��Ek� 1-�[L���A�|��Z�(`S9t:���b��A���);R_g#��$FK-�Cs��T�Lq�_��٠\M>w���[�����/���Nn�Ğ,�81d+�4x���M!� ������/�?m��~�km��ai��c�0x>\�qf?�' 5O�p��FV�R; ��˫�"��p,G`<nxx�_��J�v��&r��)3v�Ce��S0賚M��oC�4ԛ���'2�z�����˪;�ә0. =
`��"Z�.2��נ�V�җY�:m���Nݍxp��⩱3��
��a�����'��^��6F�6fJ5h D�I���KvyW��������Қlu�Q�d����8��B�����/��p1���f�ў��P�6���yd��$����"��B�hE��<Ř�!2���ey�I�� �(W/���]hH� �(43�l\Y<I��w�ax#p¨>^��h���%�ܬ������Ib�#*���4YSu���jjQ���n*?��_�u�����۲� $%׶�F㛾��U���$�l����NY\�M0�谫Z��:%��c����S�%=~'�"[d��>�&�z�I��@����C�m�뱚�p8W�{T�����x��d�^^Q�P�\<Kcc�M}k����)��(&S���|_��)fUP����^0���K�kU�OL�|�Q��������ׇ�k446&.hx~�s8����xq��E�z�#��[�3FL�E��}8
��Z����{����w��/����(��ڑ��_
s}��U\QQ;]EX�L	v�Z�U*,��γ��&���S�ƫ� ���Y_*�������@-����q��7�vh�%�<-1��a�'f��/�6��W�*յ����hX�
 ��Qp'�S@��u�&H�V6�rW��������uK-�vUW�-ǉ�6
��	�5����7��=Q7���F=@�J}��y�M���i2�-�ҳZ�9_ƽoc�f��{�~��!�6����b���J���K�G&E���F�[;+�t���� �oߦ�6���& *Te��Dx� E��I.zy ��j�_����V�=�Q��~�x���W��o��.[��<mD~.�2�q`;[zm�̾Gp��?��鏛�_�T����h����x�ҁ������A���jW!+����i���?�N�'���?����*�<d�CW��V�k5����U:�"�R��H���B�G$;�mR� 
�&��/�A&�RKz�}K�X�*j�F����*X}Jf����oQrsV�yY�Zf�U�e+�9�g#��N�g���'K�~� ��S����J�[9|Q��b����*�������N=*Jelx��'��r䯋{զ�G~���2!��[�o��BU�_��rx����UJ�HL����J�HI�V8E�}�V'�u�#U�kg}�����,��ڜ�{J�w�y���o���
E\��k������A	ۗ6�㢈:�;'��`�O�.���r��]��LY�ܻOQ��#��>���*�5�4%����獇E�������Z�hk��������\��[���ia�9�mv����К���̈�Q��	>����D�'߶S��Xb������L��W� ���1�S��3��es��*������ܕop�,����A���`��w3RsHD6�f������p���w���kU.����{�x>�}��b��{+���x�� �rOm>
��Ы
/�B�v��)�۪��dI���y��WX?���d�q�����w�U�<u�[�r4���e#UC��χQ�|*9��|�a�(q|u�I0)�0&��A$��l��U�g^��O-����O
e1ʄ�m8�CQn|/
N>u߻�f��pd䊤� �@�O.|��Q�
�	������벙(�@n����=\��u��R��n���ٵ�!�*�C>T��Ér��xE�u�S�q�r����g��&?����y҅�Z�Pȥ�#�Fã.b(�ݜ�|��}�x��
�3:�q������%�B߱�,V*�l��d<b�v=zB#��U^/�,{8�h{��ӥӒډ�R���h�:C
�z�f;P��%5}Aہ3�|�E�y*�9��h,W�����b.͆%�F^`KU�>Et�.�%(F�V)����,�j)KWl$����-�5�tE�8,�ȁ�➤`���9�ѐ�����L�f�:���u����uxJ�'6�ߥZ�F�#��M�-�����r��0�}W>.���̧�&��%���_���̅���+�$�-낫*<o\o���i48�,@t�|S�I��σM�ʤ3��[���E���]�lP�`!����<A�	}�9=��J:>��
�s79��C�~�=Xf?`L@�F�~;K�����&����y	�ܾ`�$H"5w<��+$u�4Ku�y��6b���0
�pd+9���Q�3^)�R������Y��pe�Y�߇�ag�:\�.�<�K���2OHd�M�hPlBYi;r*1G�-��eʲ{Dp�<������ h�g&�#���+,�b^@
H-tXWi'ф�=�lo�&7��˺�c�C+KG,am�;U}gSgh�o������	���*v�����m'k'�)oY��ixD�A�'��� �A4I���.k��w@���;'>�;��
�.�i��Zη&:Jt�8�T�PT����N�]�3�/� t�|�oT\I���TX%O�ta؞FWT�c�ݡK��Eؾ'׸�q�R,�i��6~ny�c ��Ӹ�+��wh)Ar��m,V�����0�{S%���k��Л��cwM~�]�2e�zh�H*Ŋ��Π��,[8]�"����� �M>�%c9
^_C�ʼRLc�!� ��2�X����C^|�4[��+�O��� ��e(mS�V��T$!����uCT��߇���äw�a���X��)���x�˿��gt���o%MM��+���H���}�T�ߑ����n���ۓ�3{#�(���mp�Ǚ/�D-��N��6&c�ъ�7��`FC���Q��ϻBz�Id��/��܇f���Hl����� [���Ï��{F�� ��u��(!B.�Yuq�:�2G�lـzS�G�6�n螸^�����Z�q'�i��Y7d��i%�$E��
��<~���nE��ͻ����i������L��U69�o�C�5�yY��|�4���)l�Z+7�݊�gOHzQ8Iz� ����-��i&@�ؾ��&����+�B�;!�	���I4�C���=�� G�R��i�=Mz��e{g�b��o"R�%�,���h��H�,u�KV߳{YȻh�� �+@ B��(���- O�����l���~Ni�ϼ�L�V��kX��igɑ~�]j~7�o��$SQ���*���to�3W$��WC�^yiC�D��;�X����RƳ��K���Z��L'f#�B�ߣN�U���-�ﶨ��,�}�
3O�`�A|�"��.\��DAϒ@�	�	@� $�HM��1���I��P��%O��L���<xG
�n{[������f���;�J�/c��¾�A���p���o�O���b���&�d��'B9�fҧ����Q�jA!��|�r��[��+g�^����}j�z��LELV��([S���6��nLk�^z�"WVs���4~n.�ȯ7�Ð�δ!;{=M_D�FDA���?�J�)��҄�JyfHR�(U�t�g������So�Cj~���/�:s38����x��;��-�����W�!����-����Y��,F�!]M�^�\��k�T���Q�{�x��N~�pd�L���P���&I�d���L
�C<=�f ����L��)7�>*��Y:�����6�[L7�N���������qHokb��	ɵ�������s�d�z�7s�9��k	Tg߆��
NF�0%j����w�wd	�ƌe��?�9ŉf�/��C�r�p�ڞ)����WI%[����V	�6
��I˪o�)@��}�@�Wwi^����#{6b�7�#�}��7'�#�Y[p]�ƆH��q���Ԕ$DLڀ�i]?�`���b�t��T��޷~}L�1��Bh׆���|��	�l}��W�h%�>\~';�P��ō�9d����S��ɷ��g�7ҞCc_;��G`�N��`�֠�}��;2����Ÿ-
� T+ 5w'�S�_���������c^�� ȶ� � �Z!���4~���!e�q+����}��O���䦮�z�;1�I�9�|�b��" �"N
��_5iN�����ʉ�_���$���/�ϗ$����gm�QU�]�d�ޞ��
��7I�))�R[E7���R��df�{����ϐ�BcA��C�.ܸz�U��k��	�`������l���cܷ�6�j��@R�D	^Ye]*i��X�h�J�d���׼u׬T)Ƹ��vq\����v+/��oa_E���U?ˀ亚E�Kg�8ok���Y48ܺ)�ֱaE�0�J=G^筻�ʌ"="e(Z��e��V�4p�xy����َd�p|��rZۼ�y�86 w~yベV��랚��i��o/.�tΞ�<͘��eSH8����8f�o��6��B��Y�J[U��s�y��V��m���첯���ͽ�;N�aPF����ji�F��t��*O�;M�Y�l�Oo���o!qY�A*����Ϩ���p?k��Kc����j�}�����<�=�����0jEV��t9��e!$�B".�'�@Di=WDe�����Hz;��7B�O��ע���R�2��>b�t5����d��^z��N��)0f�ɛ*	�No���&Ui�'#j���+B��('%P�B�8$ʌ-6[���u�k_�H������T3���մ�]P�"��u(&�V_�D,;ȭ�w��cw���;�V/ٶn
I�Bd6^V޲ߪ���G�Բ�SUX��S�F�=N
���̤CX�Q�\��$Ѳ�n`��ՙ��a�1C�"���A��M����8����
�m�1��TBzm;/����ʫ�V�e��lh�
8�ػH/��Xk�	k�9�YĠ��	+��WgBZ�����ě ,�1�mP?z&���=6���5gO~�� R9�&�5|*>{�XRΰH�#��Mb]]���<h�j#�;(���񤡭
�A��y1�-�H;I��W3�A,QG�C`���ݥ�X�g,���nu'{�(N�����ލ�i@��C<LJ�i���.䧪�RY 2;��&7m��p��g�{��jΡt��%#J��Gg���{7�-�YX�jYyͱ����:�@��f�^���s���:t����ǒ�*>榚�w v:�<ߌ�	��e۾��:#�iX^l�H�3�G���|�LI���s�Z:p��w��9�b��X��H��`�#�ub	3���&��t��m�e<�f5͐ҝ񶘵��y��߁�a�Ys���&���V�Ej^	*��^:���T�`���2�Z�uv?�^{����qX��ϐ��/��R�����{I��M��kC
&��w��!A���-5~�C�R��Uw��3k����h�d3ԍ���OM���3�ֹ�7;�����,U�jF��Ր
V8�O�3�k����ʤ��5��$2�l̺P��OTbYB//�O��� e���M�|��v��Ug�\�[j	ZrT�g|h-��F��&�A#{pU6��H���.��Va�AH/a�ʹdh@!�J��KF�T�)��� ��`u���6i�Uf
�a��}�?����SMY
�*A3,��$VJ�8�y=:ી�8!C������W�-��w=�~�}]�����W��F�P�h�g,\s�R�����c%7��}aQ3��%�.�1�&��L�_���@�a�8�O�b�-�FЗ�EmS��PP�p+lw<�� ��V���f ����ݽ�$���=-:ʕ��:��w�2���O�xY=@�	ͦXd����tĨ����N��F�����k7V]������͆(�/�b+ڶY��/�H-Tޘ�M*ò�'�3�x�g`��t�R�)f��=��4�-�|�"W}��!���0m_~���=�:#��0�t���)_�Ĺ�<T�����u�����]�e��0vw&�וּAE�┰|q&�?���z��e�y�gڬ܏t��ٸ�3�8���\`ѽzj�?G� L~�R=��v�Bn���h��������دC�|/�dn��
��
�c���~7��.�-�=g�hr�ΈjVs��������}�����<3; ȗ��N��H�9#뾞pxSu+a��ď����(f/�Li�:���tb�f�N<�F�����8�N��5+�D��i}�@�q=��O�<V>���	�_{9I���	�y�(8Wz���7�!���5(`�ܾ��d�}[�����%F�wګմˍ��n|xEf���ݣq�/�\�f��G�M�����/�sh/��I�xÜ��&K���M�� �����T*�)��m�凜�B�.-bHO�M�����L���5w�X�S`��y}-88�/x3P�w~������j��RG��ד$�6,��	}cf��wQM�J�[f��.k�@?�z��B��s̒X�֞��!Y� ���;��/��z
6�,�>��jb�,�����/��7��y��J�	�U�K"g�m�m�ԭC��v��X�����&vW�4tj-�����?�����YjRvtHB#@(��� E��|�1qt:��T��'a3��Α`s�7tdM�z��B��&Cx��3|6"S�^�aK�����l�xS�� ��L��^���"c�"E.�D�q��*ȴ�ǀ��{�15"�g8|!t%���1�Ce==�}=�k*�1����֥�Z�cJ�"�1:H����F�jLN��`i"�d�>g^�Q��
�݅����@�j3/��7"r'0�$�Gme�}��fgE�:���)�f���L5�l�1����N�H� M5��I	OSέ�F/�Z�[�����aO-�''�5�����N|�vb�����0��p��l����<�G�2��W��m]s�����s���1.1�\t/T`*2���������:l*Q�l�[u,ƨ�X�aw���O�aw�-��	w2$"�u��2(�����xe_c�y��I
�}��*ߵ��JW5ʯ �Q?����i#E*l�3%sR�A���8�I�ch�ޫ�B7�T�ɷ��SS���M`�a����-�}���x��$z����Jl��N��E�%��k����n��4]�mbD�
��q.�j�} ge�#�s
������ma��`��x���^Q"��^*�SƑےdđi��Ū�K@��	c2Q���i�n��X��ojs7�	����dV|"��ؖ�c��jr;�u�u	ƫ'�O�#���:#�������l���������T��ݚ-%{��n����+�f�y��V����^�;�Ae[�4����e��f=��p�<��?��ʴ!�;�mʦ��r��W��3V�d�pD]>�^�D~����/1�%�U�j��ܮ��AYK����J���S<b
¾H�)�W2˙U��~g�㏝q�!+Vb�x����l�;��2uP�h�9�O���#�!�H6��G�o�`S�a��u�%g
8wN�V���<p��A�o�cj�5t�r�@�.ØC��G;�C?}Q���g��!�9i�^i�" o�8)GL��&�A��4�M�U��J)l������wʉ�JZ�Y�à�����b5�e�;��DK��8�/m�`19�F֕�pT�JW��I�mp�'�*�H����囬��Z����cZ�:+·w�d���K#ґ��=]�Rֽ���ux���;������_7����56��4��@���������F�r��P�zp���`��0��ff3B��v�{s��D�����s��R̵z�Dwma�&4�Ǌ&k��j5�"��~���$��h�k5D�B����V�d�Y�F,�_��P �q����;�+ݟ,ÃPH��p�q� ���[�& }-|[��=On�q�#���ڌ�����i�����,��Ӑ�3����aH+�o�6˄�h���.2'bW)-�]ٌ�y36�vO�yf�Y�$��x́mxE��t��K���p����1=���O��z�!�4�>Q�@ s��\�E��"?��`h;�uE����e�÷���jV�ԲC䮷��ڻ�][���t׫��\��}��E#�Q�k�EJE ���GںF���e� !�i=��MAnO$�a��y���򫻥]�§���� ͜���O`�%�i���{�+R]<7<��b��{��js�D�X�:��� rN��him���"�����c\�cz��������v������L)�w�F�A�J�Y7��&@�۾�5�p��jGV�$�u�W��1-}z�ɍbU)=/���'��,_�����	���w�U�;���o�L;*���;H�씚5G~��g#��1�`�e.�S�߀d�ETgλ�������K"��C�� 9@�����E�kXZ���Ǜ� ��g6���BT���D	_��< �(�.mI�/N-���u�_�:D���ŕW�y쏄��K1=�����vj�����v8�Y"��tk�:q�s���_�E�ϧ��6^�[x�ӜpL��N�P9��=D���!K���Ƽ�h���3��!�JQߣ�����O����Ւ�(L��.pҢ9x{[�o�Bطo�X�6e���<k�u
[K��X�"��B��4���ؔF�\.C����^(Ť�qi8:y�?l~Y����H�\���Cs����-��������p�{���+2�.�,,*9$čy�\_�^B�q�K�`e2��=����a�=�ИH�P���L��B���7%m��Ƅ�6,ej¼h��Ü��By�/��l���G��"�T���F���D��(M+�e�eY�����ՙ]b�C`��������Y9i�B5>p��F����O�OZ�� ��ҟ��eFՌ�H�z�J���>�d����8���.O-;�<,�c���j٦Й��7Op��;���%��ҿ>�a��@r>��Ɗ���ɛ�p�6鯥�Yf����5T��hcϖ�˴L��z�m��c�+X[7ʗ#R��Jc��o��B �3
�`�Nxr7���ۘ��5�'ռ2�(���vm�0�q�u^�
��l�	C�v�ö�jr(��$�)�=Al�&�h�!=���hB�EѺ�GZ�PL�O1��J��	�Wo�e�h3�F��ɉM·"�{r��1�߮�-�b:��l~��d�gC�z����N�S�f�U�4�hWs�g2����V�^ cbU"�$m�u}z]�Q5����O��"��T�l$E�1Ģ��h�M�e���$���K�'���O����|l�����6�}1������_����՚�?�}��?�h��^��e�v�"���s��E�X��	l=9��<5�<�!x���g9������t5ٶE����2S^Z8��=�u���$�EMi	خECN�J���$r�r�E��o�nRR��6�55�5���0FZxw:$��A9APؙ�h�;Sн}�ˮ
=i�hH��;ZiBr��B#w(�����N�ҴCW���@s�jh��
�,F��,�]�IW"��>�m- 2���Ah� �!��Zb�OoN��8:�(إeŒ��3�h���y�>��ȯZ�~'���5�Z�!� 
�K�ad	b�5�����Xz���9��_�Y���`�m�m�+t��{�A�����-��E�ec�ï�x���5�����&�LF���K���R�B9�g�ŀ�G}�0�3��l��$J����Iu�g܍���5�9 �2N[��qg^K�K3vk	g)�����r��P�=@j\��7z&�o4|��x�B�	.����N�2Jr�
m[@��� 8���b5�JȨ�O�O��)�Ⱦ�/�a;wP,S�Ӄ�3�r�G��J����*WЄ����u�7;G2�g�������]qOs*))t+��وJ+qG2N>A������>e�Ku_��$�@�:�Xo�4�caV��S�C����H.�
2�4��%<���4ⵏ�;d��
�N�rt���d�ȵj�3�ū��R��1f=1꺒6�K��-;d{�L��9Ր1�=}G`����>\.��'qg�������k":]�b�|�l�g�`�n��˖��*n�x���c3��߽8=ל��w!���'�L�yj���t�n~��*y�x����q�sdA1��m����k0�WH�!RE�V��Ň�e�y
iv(Fg�G>F��1�M������0K]��jΛ`�*/EҨ{�:�.%�����}B��Z�*���,��ć�Ƶ�!;S��� k��'�����������]V{�mLD2#A���=�����A�E��T
?��Ҩ�T�1��6�M����p^���:��#�u���g+a�#B�c�0ݮ�3��H���QF�	�n�V@�v b�:�ޱ(���n2�!�e�#+zb�����g��PY�(E8ﶸ�q �Vcm5�>m�rkGd��ky�ĝ��0ȼ�D6�������|1�mnB�l�8E:,�~����7�7����j�n��
�� �bJ�<,���f� �����X ^���Ok�)�Kc��q�Nit��tj��J����B����N�dgT.J-W�\Q������m�|�'���M�QƖ��I6G�=t����g 5�E�K(6�Hf�~w5�5�J�`.�(t�}��\gC��=��s3�<���v���=-�㰊b����@���ܲ)�{Z��� �M��%i(������z)KX~Z��`�.����;^��ND����祖o?cˋ��S���1�~�;S>�������9|-/pr�2�Ѝ06|_異S���C1p�y�Z��?�uN���_p�e��xJ����M�',�l̥����l&U��p"�f,/]t��l���s�N�:h�j�ac���������-�I3��__�MS�#�'P�A�p�v KuƖ7[��`���j�m�wg�_�$A��Vv`0�@�:S�����i+�L�?f�w��y����+b�lm���r��@t������\��&(Z���yZpךmj��L���y�׉Q��k�4kY��Z���`~��Qv�ǦR|��Uªb�%) j�B������~K��<0ž�ڙ���Z�e2p/����*'����#����޶�C`��'�]ע�e
Qr�:jjHc�Ri���� �U~."׶	�Ḙ��~ �(�J��`0f\�ǿ[X��@���ӣ����X!&���F�j��}�{�d��ڑ#�jrm�h��!�"k��W�Tݒ=:p��a���_��zt����T�Ө�<�HY���>����͠�-�h���o����[rw������紪$T�ȭ=�[����]�y��f"R�e��2��u�}f' ~�iLYJ��i�ڝq�����ܑ��)u�R�g����Z�?��F1;
ww��|a'������A ~��fY�������J�"yg{��~8�M6��.���y�c�_J�����ï�s8����[@F�\�$-I�L	���z���������sr����Oկ�<�8~���U�*�ߡ�>�M�do}�s����%	�d�7W�>�N<,|�Pw!�9Sj�ke,����)m�U�n���[�����M��%WfV�?���O�grR�G�{��}�م�������ezs���T��3����g^�?K}�ѡS��z�Q���x�-����r~�?T�z������{�9�5G�їV�q�2P�-A0���y�Qf���t�,[�,�aZ�QV�U���E�~����g�6��<�		 �̫�����~Y�I��`�t'�\m�d�HH�洡�"eǵ�|������^6%N�%|ZqeM)�%�V����x�j$���̷�0��";�yĉ��ir��h����K�U2��l%��h7IM>����5�僦5͜��0RGy���o�'�
��������cz%���
�f���)��
�@K@YD&s�;�B����:'@YG�]��آ3%���2��a��o-��(�}68�LI����kZr��}�P;��L�{c=���D4���6E�*5�p`�ɝ<�1�``�*`�b�����ج6d���D��[�,ԁ�Bm�y�ȓ/x�����׎G )�
��x����j�h��23��ќհ�Z-f����Nv��'oߍB]�FD.�e�yH��Y�K�PI\���GS�H1�pU�] A2�u�wG�CUay��*� m�vW�b��h����LIL��]b Qj�Nk��%=7��F���� �\T��O%����wj�]��f�w>�ɝ)�@z�(���h��l�i�)<��?��4\�(
�N�����S�C����15�Rc^nVo��2���M������>U�����vW���}�0����o��{F����*V����_Q}�u�͉�̻\��8��;<���z�̳���gM�;���ɄTY �&��o�9\��}
����%R��	���<�~�#l��Ҥ5
}�>�Z�L� $o�l}�A�gLGJ���d�p� h�2 ��
9z�И���Y�����3�a����B-lX�4������>.֢1���ε��Pdc���2����:���Blz��6iwh��z6�jŴ����6Ə�ݿruj��W}�칱�Eo�����A]�Mo�TeYo{�U��C�SHʮ����*7	f%��N�LCL��/
��i���i:ain;��JT�n3+c�N�s`+����x<�����!jJ(+S��5S�
,������ tW�t.�C�*�ϙ�{��YOƅ��c�G�K�,'QI�Q��&.����
�[�e���aG����v(�d3cѾ��m��?�0m8D�e��`� q(�vLv�9��f�4��h��4�CV�[s��fˇ�uZ�xc�3�����a�ε��pw�����B�H�.�8�u��)�*�#�aC�'�puJ}�Y�7×D�9ʍΞm@Ύ?$�i���m�+�+�3z�cK��7��ˊ��$J��e���~~���0�;h��.?eu���")���I���҄$����	�㫜���n۾����:�jS�dR�WhvM�Zv|��>@㧀�'���r����^Tn��F���jO�1���Z_ޟ�P^��^m���}�����\�)Y/��(j=��t%#�7Nߋo�o�2{�>��]��G��qc� aI�m���6<��5z�C�S�
�qG��}]���'�⡜.�b�1���p�?>]g��H�e�`B����D++�B |�;h��5�j6=�	*p�%Kr�	62pD�ٜ����G-ޡu�3t���K�}��S=�xV��tJP���^Cj��w��_$�+�wwȖm{�����ᮃm�V��>8}Oڅ�a�*_�l�r�h��c��+�K�'�K�R/���\�1s�n=������+F����+�Z?�c߈����6}r=�)�6 {�|���1�£/%t���D
 ���MF��MGe�N�[��J'aCr$Ey.TbmD�b�&�gp���i�2J��E]� �c�`LZ��R9�}�og�b�稷�18);~l9W�����ˡ��=q+J#;\{�2��^��o�|�6�U�����
xn�S�P?oHf08�n���0̙oPh�[�a7�^~V?n:~/�￡�5�u@�ӗC�'�'� y?����q8H���iHX����pI>��P �B�"��yk}�c� ��yi��{�H�k4�\l������(30�	�(e�	�h<��Ŷ��&�Pû�S�e[v
�|�e�_�?$�r����w��^�Z��ס�v���g�G��(fɹ��`>��de���H���gP�*^Ə��4�d��Kw����-7*%����ƈ ��a/ؿ� �|>��\S�"��^��ĥڳ3ݏ;ОMD��E��Kw�z��}��Upy�O9�{}t�_�iGT�rZ����Z�j�m,=Z�;T�=�:c��f���������֧�,�?���U��m���g�q��Z�ܿ���@M��o���~�bk޼e�6���%��o~��M���fC���΅$E@�4|c���h��6�)��eSL�I�@ m���Ф�)�������L:�R�M3Gd�jwu�x}����=nY���$����(��ga����bE���L�|��(.
��_���!�8qU��x'[=R\ȉ���Q�FQ���iS"!_ ��}wmx~�����z��I�΁��!N�CHˆ�}&��TƩ	FԪ5����P�IŴGm3Քۻ#q�����)HҸ`�t�M��{�R}Y��J��yǗ�k�W�eW�.�eRL�����M���pv;�Q�w����!�_�2�"��(᫪�%��v�.-_
'��bBg��;��An�i�iExt�g�;��#��2CC�s��^`I�ݖ͹�˷>\���8[�Kߪ)JD	\�j���b5��l��[y';���i������0��I�Q��-N�����"&a$�ft��6�]m1b��W $�E�qٝ$E�9Om�mJ"��9L��k����儊Z����vu��T���
h���To�$i�:yHJ֋A�jP�&�o���"�-��+Qsv~��ߧZ�����S�]-[_"�P��N-3 ֑�y���>*��w�J��y&w~�ݞ0�/җ-ġ�)l�X(r�Fm��,I��g�z	~��X�C��b��*��l�с�E��0&�bq"�Z�){�<3��[y�sɟƷz�{z?��~�7c�����>�SHNz�vg��p�|�����e=���W���א�wUϻ�ƞ~���^v�{��%~[(6�mx���:��qp��T������c�Y��Af%۱�CiXQ����c&�>�cա2�8F:"�:2��TV��������������~>�e��FH��Ymt�:��S�0F扖5?{$��7���6�0S �g�TE�W�v�ZT�ຝyù�(����ki�'Hc�U!Q;���I��)�r�9G6�cR~<�9���)0�[�3=�)N���j;^����\L�^2�n�x]j�ՠ�_�G*A�sg(�·s�V�<#��ie�e5�µ���7����)t�y**���l�t+q������b0D�jB� �E6�{K�I��|����,��jɦX��;�L�]v�M�P)�~Y\
1OΘ�~��)��n@xȽ/tR؞�3�H�.�Н"	����;��ęF�@�ʆ����(�Y�ڮ�c+J(u�L2)\�9)h����w#@�,9W��gs�7����|bE˟�(,��B���0⠂�3%mE��|l=:��|��,�̥�h��tI(4�%����@WQ�T��%���G���Æ���!\�ɎA]����������M����`18�k�"��)bcEJr/����+���׵���ҞO��1�5AlC���/4;hL9��/�WPw�b�t¤��@D����c��Q:ek�&�R��E���7�;[��T�[S ���k�}��+Q�E���w�娹������r��U�e'4�ʼg�9���6���Y��&�k�,|q�D�־���Tj�'i����*�݅���'O�f>خ�B�~��#���b[):\!c��E� G( &��Z!�L(��Nf�@<Aȕ�l��-�S�=��j�d��v��-$��	R��^~�[2[�8��3s~�|ŝ2I�#Wh�X��NP#C�{S��~���=EJ�\{d��:h���I��Df��� ��n��J�;�
N�9��J�z�vQ���;����c��(l�O���L�8����%D"Dt��ٕP����P¤�V�M����#���~�<K����U��w����R�`5�3R�#m�X`�O������'����'e/�8��I���AC���y�2����[3)�����o��d�=�4�LY8gC�����2ķ����~��b�ː�	��>��&��F�������O��n�|��v����zhce\Z�� <8��'Q�YuG�a+��x���w<E���uR�� uf؀���$-k[\u�0r%�Z@�v��&i���93 ��^�n�����z�%5{�3_�  t]�D����3պ��|^Z�a��r?G�x��ĽV���ܚ9��c@Rh9L _X����ݰ%/���;s�Ђ���K}��Pq�S������[��Rf4�&Wњ6�I��}���-�����5�.P8�;���eqU˅��K���~����j�9����s�'�P�d�%�Zt�c�@i���p���iJ����~O�w|r:��u�ࣸ�Mw���p��z�,J'�6F ��-���:��s������E{�e������9��L���/Jn}O~����f�y��~�o�P�������U]�s?�����G�Oe���Oj���r��/^�#�Y�I3@�( ޚV&NW�h�����vx�+� ��r#����� ���x���d"F��9(-z��.�;2���]��o�t����,��k^�U���Z�e���NG�yՄ���~�w��-���HI�V�UXoC'��L���|����d���s�`Dz���I4�T����3z+���"��3
U��gȁ���d��ݦ�Ju��L�(/�4f��:�	�������2��TG/풔�7A�
Q; !^��W[����lĝ����as]�ُ.������=�7Ԕ�=ԯ.K�2�&����ZhW>�M�A�m�藃1j�U<�C�)�:�9�%y���[�G�|�ˉU�v�K[�e�M��'��.@�H�&��ɲ�l2�+9����&�;���DB?K�4�����2y+�Vgűs������)r�P�Z̹Ç��!��
Rw_W�b�F���/b	
k��0)a��VH"� ��������+5s�<uLL�S|�6�4S�.QBҥ{2�����B�̤K`������`Y�Suf4�^ܓꧭ!?��@����/�0��ù�����O?j�G�Y]C};�����J��T�g)�%��8�XDe����Jv Ԣ�Z�F]��0����U_�����)���A�+K�{�ٿw�~��+jw=��������N��oB`zo~?p}��������g�߰���/�A����e}���|!��9���ͯ���ܟ¿t5=/຺gQz��e��E/��jʪ](��+�=��«6�m�:q�
�D����r��U*~<�ɞ3a����`�b]����$�O��!����;l����o=��2��MGe詴���t�}5i���&A�,f�\��?�FU^:{~W02�6���+	F%-����űi$Ɗ�֙Żv:
sJM���g�X�P���zG���싔gG[���j�N��Io�B�@��TgZEM�}�{{hrP��#�MED"��G��ټ'.2�{w��!�8�y���@���h��Ea�u��ӟ�kDQn>��V�Iy�͖G �R�K�R3L�iu�[T2ߜY�����֯�&��ϐ�b��H�S�5�~[�^+	<1bC��s�]F�w�flJ�S���:�  d��L`?!����at]��z�p}t_Y��`����X��+�:�M�b�`L1R�^�h�d�;�צN����]���9l�TdC�U��V�=�;Rg�:NjW[l~\�wܹ�����E]�3n�m�?���|�
 �힨�bjX4Ui�-��S�ƌ}[���t�=��i���.��ز)���)�LDЁ�)��h���gi����c�.�Z�4�l)�~g���m���Ip%4�ܺ�����A@G�^[�ri.c�����o�1�	"�h�W�}��*���r<�2���jg�u%�1�C��9T;n�/��g`rh�d���\U}֪:�ì(����nR��9��f�Ņ��{�5���6�6d�N?l��qol]��������L���'kk��L֝�w-4��]�=�����X.˃�ޢ���1�E��ң�LUH s��/�Sw���xȌ;�R
��y�aAI��!/R;����,�ea��g>aC�D����ښ�%f#;@&��;2I1/�;t�=�����l�y���P9<E��x��&�CN��5�Cf��%0�g�����ӲSK>1��|N���Y��)X�#�T%_ߛ`� ։Jʾ�P~Jq���ժ��`�7ٽ�t�-�Hh*���Q�D�<� 򒍗��hG�0&��VZAC(|#��"�ׅ f�bv��3��s�X-����Y����ɩ���5��7>4�6�X��^��C���N��W"��
E2}�A���J��Y=X�[�>��g.�b�^�*n� �\�=���&x��(a����������ZVf��@,BB�P#�ֲ����õ��Ň%�1T{�,D"����"� ��+D�76����&�PLw8��F�}	&8ϴ#!Ac1��B�?V��Z�"�x�+����߫ȿ�&�����7t�'� �}U��嵋��� 7zϹ�eh�(n藜T�U��ʦ���w	6�Ab�赐��\%Љ]�������GK����%�Ps~9��)��%�J��sfda�؉Ͱ\/ �r�����Z�I5O���vQ���ʾ{&`� ��c!#]����L�76�:���F��n���$l�):����~Shi��I{r�$���G��y;�c�=b�w\Y=�*�O��|_ZKD��WI�<<wC��V1{�z��7��F���tG#N���#4��݁d+&�Heݮ>�ш�@�P+���4g ���I���	�@��lO2A;C���I�et�ܥL���F��m���E���_���A�_/A26�q��M��Jh��� ��I�/e�@�6���.�1R�KZ�4�U����e~���Q����jv�¡o4b�)��3";���8G8^���]�g,� �5��5�^�Xm�TO���jjUxȼs�ҋ ~ccw�:����v���$��E�OR"2ܝ���;��r�V��ƪ���\p8���q gd-G��.&�l��y�L�~\�۞�����xF!�c�����F;^�!rld/�R������PGȨ~����)6�`�8��+��v��;m1��v�"\ D����=(��A9�qYQ�"�7���95ړ3�l{�\ߏZ�)�b�gl�֯�[7�9��H��DSe�L���2�V�uO�7���q�*�����B���fB�/��^�Np��( ��rlq�vG�,c��L��G�_����+2V�/:.Ԕ�m�ZȊ�(�0w��o����X{����[�$QEl=���T��� �����K�s^5fH�i�qQ���]Jl�ݣħ��sD��ʍ*��V��E�ool|/��u�Ӓ+rU�K��LS�Ι�N�*�~�Q�7B ���1����.oXP����G�T�%R�h�b�;V��<�N�j���ꁒ��ͩ�!׶��O���+��}�;�y��~�tk�*9�s���f��K����������r=�e�Pr� pVFyu�|꜁$���|�9��N�qHf-�U@0���p<]��,�hj���W�[T������6���HG�$&5� Y�Q�`y`��G�.B&+�.1Aj��d�w��OL�z�sW��ў�I��c�d�������q���!f7%7�����WK��LB..zM-e�hQ�*j�
K�k}`4��[��
G���#�Z��I�|y~�t��[ �"̱����mFD�ә��m��3ւ�����\z���9�1��G���7N�FiS�Hj	�k�03K�uEĐ%@(����>w���$�|��=��yΟUk���k ����C�:���+�!+�A��&����JAh�����U������T��+�y�;�y��<�F�7!pf����}��GK�.�*$�$�|F�a��ߤ�P���*���Z��-
�s]��6[֦��Ռ���� W�BTefۗ0�-��C}��4U0�����E�A�d��3T{y�GA��܅����Q#���]�Wz�dǵ��
+����E~*`�L>�q���n�u���A�#�w��԰+r�b�Ԃ����r�����C�Tx���@���υ���0��g_ٻ��I*v�<r;�$/�xiM�D.6���R�!]6�x�'��6�^[<���75�4�9-�F�g�&��x)%�oB�4ߏӔ�{�W����ѶC{r��%/�,���9Zݧ|q��z�P�b�,�*T���G��)769�~�l�ޚΙ�][��q`s�����������j���.5�D4��%E*t�U��d>����U۩P㫟�5�
���K9�=���P�Y���L {a�9�����	R��[C��28o~���}�|�Q;%�5�giC�`�aS[\���`��%KN>ޚ�ٟ�3��*&�4�l�4g�,O�����yt�Y�5�
��k������eh�**�f.U�I�NgDr7�	��H}�$����p{�����\�w 9��k�����$\`�/����n*2y��&��2��3c#��|rC7T�\���~��}J)Y$˰Y4�E�󣜤�����;�X'�삀4��`jVD(L�9��o�0w��`��Ɏ^�Bh���#����L�D�p��_��~]���/כ���'yy�5�:�|>O�	��!�����_e�69i�KS���#r�g�C������?$`�#��t���қ�1}���*RSe�~mp���M�#Esk�RG�&l��F�Ro�r��V=��4T?���f��Fس5���<�|�99�ؚ�_�0�D�D�����@��,�K3�����c%y����z���T(�����N37K�H`T���v4-;�s���_`�Eɍ��|��ve�2r�3>�iA5x��k�a�.k�n~*���A+c���+1%)Xfg`
+�'�ezm��ȩ���}�N�{��z[�m���T���,v*xa-{�Hn���d�ۗ!�>+:>8�si��L�Wu�����y1������s����
�ue�6��t�W����$~�������k�|t��~8��C��jH���D7D��ay��sٺb�R�+���S�T^��&�{Q`�����^��Ùx���'sq4�8vX����m�2�d��EG�����id0��@����`������O�� @r����;Z�H�6�eN���7Tf�����j,���Tsi�)�Ӑjؼ�9w��}>B+�r��@~�4�ؓ�9�7Yb��4v�s9�������_�c��-�-�`���tI�q���cUeI$��(Cy+UoPʔf� N͘��A�F�.�����\�T����d�t�Kr(��~�C�����.A!fN�h�-5�B՘$�?����GrX萙�Ö�UKp���� �@��p��22���,�W�|���q�Y�P,v_��lP�\#�T�Z)X�栋��Ͼn,�����R1>e���9��s � |Da[�R����u�����ƅ���Ti�Չ|`cƢ�\�6-y%���(��8N��DЮ��[�b��A����@�"��h q�� u=�Nz�]J
����	c�x8
�]���c�(֐��IKP�s����Of2{}�v�#�BQ�r!-�U�XO��s�x�<7E���m�R=�_���2�>�g{��D(*As(�/3f4�!�d��K~|�˽��ǰ����7Z���9(º
�����Z��8R����^֢��Nj�U)�:xP=fYmhtHrnn!;���?��u��q��vi����a�ډ���
�������7�M���5�7��/�����H��x�h���pa�д��~���� �n'�@6:ր�����|A!���bX���L����z�A�M2(�Pu.S��c������Y��)eӦ��?"���pL%�q{������������:�1~<ڒ�#�;�G&CH!"2Ȣރ�� ٦7+Y��ҫ6˽�{��m���dӆi��<�Q��
�d�%� ؘu��U��q1cP()b�@��!Ǆ���R��s�w&����e�̻9�X88�M��jX�)��i����#2�K�+_����[p�~�</r�BS�:���1&���<&�a�HDx\Qd�[|&	�T�5�����7�5�FaA�S0,�$�)�D����-[`�vd*��L����"zYK�kTӢ�r��(&Z�YD��gצnK�=�CQ�"�B��@�j��;W{�I7����r�z�h���	�y��ʇ�Y!���Ȋ�Jy�og�>��gex�ð�����z�d����Ə�<;�Э9N)|�C���n��U��~�6���If�A	�p�>w��\�T��u�����L�ߣ
�M�i�� �)��XJYA�Ǿ��1{����}S��D���7V��$� s��!	�k����X7Vd�!Ȣ��jtSr��Ϯ�sX��m���;�x�,{��T���,����{�5
�yy����u���b�Ŵ���t��*TN���K�~U�I
;�65��?1���<�2��g�a�5�eƳ���o���F���gx�$NJf�4����p"J`a�
�NTPWy����{-����(?w�`���j��w��PP��Z��~b�'�k +��O(E�9�!@ooi+W$�9��t>W���<	�"��M�p��*NQ|Cy_
�B�(��8�
��U,Y��r�@-}�~ZDa*��¶O~cT�]Stڤ�MzpuU�?�ktB�L��w��x��Ò��rz����+S�+f 6�]�y�����'���6V�X��ΏwcW�)�
M�4�L�T���ǖog�2�{e��V��	s��%=�<��2	焑SЬ�(1���w=]���e&���Ga��a����We%$@m�ю5)A��H�9er-�G�guR .]I�ku�	OM�b� ?^�jN��Q�4�8 3���� Ǻ�.�e�p�o�-�u3�N��,�o�Pw�(���d���#��1�M���e<C"vA�E��K���}��D[�ǀU`�Q���c��~tQ�,z~Bط|����#��+���ʵ�$
�>)�yze��C/��;YZ#�k�����̿���|�&fk.�nr1��7g�����Փ�ޫ8��P�'��E:^�ա֎���1�l�FrO�X�ŀ�Uc����CvY�W;�y�9ر�|S4� 6�ž�>{y�^�{��q�Y�$)�mN:f�{���W�U��/I�d:z?�+G���\Y��}������F���}�~x���C��o�n�)o�닙����u3��;��"y�~2���B߽�q�|A�V_*,���b� �D3Y�� ��D���@��J�}���i�e#�T�P���k���m+QZ�v���.�X�,L�,]*�h1`3�����U��r��j�M_+���
E�S�]eO����[k�5���$u�a	��
J��M������ϫ5Aq�z}w�i�-S�3�B�׍�\v�5�,�9$oߵ�_�U	�}&
�	Q��h6J,�f��Hm0p��2fW��K i{��Ac��el�H�g����gݚ��Y��,��x��Ma���u]3��pF�aw������]��]��� H,`c�DE��T��L�j���_������xw�ѝ�˥����^��$xTl�_��CRҋ`5��vt�)H���������4���6f$	�'
�=��W��d��y	�R������Hl9�@g%�R�����[NdA�Wd�ŬW��������A�\�]&����~Qn9��_f�4$�.��#;�����ޭ�}k��M�������X��4�񿝎��WL�+M��9T���#+ě������ˎ.{��f:z�h�X��
X�&��5_�ub�?a�V�os�ㄠ���<�����e� 3�EӁX��"L?���%�;y�~�̜�ز�+tZ.����`O�UL>�H�
�����-�<%F�t:�^~B����~�����Q�U���o�<e��ˏ��Ζ<�3����g&9��詖G���F﬿��3���0Y'��vlY����KV}���'�F�F��1�H�k+�lA8�m<0��$��e��5��ˀ��FZ�����(TC%�f���)�r�o��h���"��s.H����G}_؏���~�B��#Ã%.@O��~��3�sI�� ���<�<�o=;����_�9M<�$�]������� ��9��#����u���֥P^=�G�\�K���ެ�M�6��F�c7�)UL{��zK�
rS1�օ��o�H�QQ�7���E�7:�۟�й��B���
��,K�`-,bLlΌ~��F9�V����yQU��`�4J	��� F�=��'�;��X<�ғ](,�L0�K`�rn�}OJ(s4��7���*�^#`�����	}�0/��vYi%l�H�[��,�4�8s�\��%��Zy)�N�*>��_�M�6���n	�D�����|�X�� �7�J��W�~t7vv2~�Ku�����&�@8�06�7�x�y2L_�����N��B5:Ԝ�r����Sr�r��#'aa �"�@l�kc�o�jL#��$�qg����_�I��@�tx�z�ێ�kR���`ʈ�"�>�Z-�&
��k$e�XV�y�>����|��R(�����`��z�5F��"�@��|4E��!K��
*��^��xt�#�_JP��=�x	��1O�����/r�!ǂ,���sz��D�-�of�թ3�~�l��˄{!$$D5p��3���o}:�s4���9[�Xf߯��T����ˤ��\�2�^o���,�Y���p�k?���:.�)����.�ɋ�tf���3��tD}�uEj�C��T�E���=�hg#xA�e	f�L�z��"]�r͆4t7q�!]��^m18{�S��b赤�l�s�B`;�kङ��\���s�Q�%7{K��-�����͊�@2��HW	�#A9{ ��n�_�����q03�&m��0o��>!a���U���7���Psd�g۹�,E�g�=@�o�J�C�	-��~�$lB�*7%�T�4��g�#ܫB�Pa�.�����=T2?��@�sTǱ\��(^���%��4@�"����*�^�2� k�Uo���H� A�����}p5&;4UX���L�;:��2u��| M�U�q�6r���|ls8����k�_)&�a��+{�t󧄈�sĂ���Q�8=������v�ǔ�*�0�=h1Z�wU�L4�UqM��愕f��*�������Ή�o����@P�
hc��!O�I��866��Q��?fv��37��V�gxa��%q�J��[{�æ@����;���	�ڌ��Ɓ�~�F�I)~~�����@����z��71T7Y4S]���*��:��;Ι9��H�a,�_��:�j���A��<�ʮ�ќ��_��tΏg0B�M�39ՠ:����|���.��������R./��1~�կ����;*�XR$���>Iw��쟨2VP��_;���}��8P����hw�}��S�^����Z���(�\l�;^�W|ؽ)4�(����	�%����{�kO͕��@�O��$c�T���qM��9�";S��̉��S�[]/�_��'�Gt���8q�'P��c�=��z!l�R�;R�w`h���l�a���D��H�8�֦���t�ې��g���;�3_Cv�d��U �
Dғ����oJb�����I$g�=iO�A�\P�A�X��lۤ׆��P����Qu����0��l��h�L�Ӎ��IN�t�lY�'����h.^�K 0�
��fe��j4�����)� p�ᴇ�}�N����F���/$r�ty��}��9�e�F��ɎB��Ќ�����;q��]��׸��I�T1��N�ߑ�խӦt��)�,��CJ:Hx�f����x���ơ�!G���3S4Ծj�5!k�P�1�̩�|Ea�� gg�:�D:��B�&-ߒ�^��ٻ��愫1.qd�7&4{���@]�~�P��,�DUFH�U��8�D��Ԝ�����X�n�:u摎�1��՛%��?Q��KyЧO
�!zpt=H����*`4�8ء�w��B8�Xy�c#H����'��hQ9��z�$Q�����0�
�\#�Rw������.�:g��~��f���Z��$�W��ag`�<���'%��u�j�>�0p�
-��&��ǝ��ߌ��\�Jl�Ѹ�w�n�@��%�0�r{�=X�"��Ze6y��5O�e����Ƽ��*�N$��=7������h( �mpW����/J�:M]�9
#� ����)�c�BMU�����g���S��������S��>|�^��6���ݯ�h�r�7�E���~��\�sS<��;f_���V%�J�0�.ƣ1�X"��� .2�'�@Rh� "cK���=j���[&�o�VZ��՞�%��%�}ˑz�D��`����M%CL�L:βu�[��s� ����Hq���۷W�Z�S��Ѿ��W�8
$ݵ�o�0�
ܼH�[���<����j����w@pR�u�[.��isgo��_9>A��Nl��J
S��/嵲�]w�*cCg$AZ'�j$<O3��ɐ���{O�EEr�P��g.��A�i� ⬳���5�0�m��:�1�s��]�M�,�$�g�Ge��Tt����Bz@Ǆ���s�I��3��vk��砓��Q����'
�X#��4����m�4~�a�\/�@�K���r�v�q�vY/CN��rj�a���*�y;5 q�	M�2�&h�5��D(@e�����M���$�#���/l�H|��Ԃ����'�V[xPA"�d�������H���܊9̈́�KcL|8�G[�Fݟ���kr�pD>2��d#}u�'�*�E�ɏ�)VB�ɟN�5��F��c1���%�cWs4`��#r�yoQ�����򂨅s���U
)�H����ft�҄{�+v�'�9��4o�����J�M��c*#��_�)�B4(�')+��#���d�.AP!�t��5W�jH�9�U��H �K6����m�6�9+��k3�3X�=�n����wB���/QnNي����SoY��>�y�2��8/h�4���YQ�D����I�����bm�_5�~�w���F��k1�W�l��^��qZk�)�5���X�اV�a�vpO���f��y�> 0e�%\�hҏ' �WӾN�e4$�hS���K�Q��lde���Y}u{̕6)��G��{_j�z�k�M����,�� ��w&"��y@��mzatNo;���2_�u�4T��X�B�.��=wI"l���A��1�[�J�K����j���EO����ːe�"9|��4 :���������ݹ5'2�J����c8�-s�%ɷ�64��p=������ˡ�	ħ�02"zS7�g���A�I���'�+H���	O�x��s���<�ד"�k®H8��{�XEg�v����O*,ǆ4����Rsi_�p=�;��C�6�5���W:zF�M����ݱ�)52'�'_��?��⼳�L�l�,$�a�U@��.�����{�Y��HF�$�w;�Udl��-_w���Ki�<
�>oӶ��} �5ܨ~����߽-
�<��Z޲�1wKܯުur@)�q�����u���ո}P�78{{�w�p�cd�'F����c�d��L�ڏ����:�j��x.�Y���vр�����
�U�+�aG�&�I�g�*�ST�=����6W�|������J�^�Q�W�WhG�y�e��ۡ��p�!<�#;V�WZǿ���2<^]�Ȳ��x���R��P:�[k�:����O��h�M?7� �)���
Ư�l�W�6��߸>����76����z̦8h�H(�c,;�v�|8���#�"��Ⱟ2[e�H�t��N�{�W�ք1��(��s�x���OB�ila�1�ˤX;�)A�B�<�t��r��1�|b�����q ٞ�^��s�F���"gk�2�;�$v�L�&Q�@b."csy��V�w,Y�1tv�k�X5;�i���k����wAh�H?R�_�۰�3���9��r�z$|h��c����s��7��P_��j�#'�rp���w_<�w@z�&�
�HI{��^M�zm�D�f�.�bx,Q��'�D�i�Ia���x����S0�!y�A�����NN� �c
_<����r�r%�n�#�(�g{�s�i���Mx� ��eƊ�HfZ횭o�M><Fj�Í�H]����C����E�Y�F� H�w�O��������G�r]񩙟s� �&�����q�UWi�%�6+���X�-tGO`N}kp��y�r���}����yw�cd���>5�mb���	��#�$<g�c@�5�Xy��+t��'�0�Q[!�Z@aQ��%�L�8��k�ݷ�\���?^c�mޠə����&���7�áj�;9�I����'k�M::�X�MSC�����U�^;p�gK�.G�F�;Gx��y˧�@p�(��R
j����2�1[O����%*T�l�������Y������5(�/�}�4m,���HFo�\~�!�\�&�[�TcT�Wu�W	^��2����|{^��~5�q�`�qQђ�s��\�T�rZ�g�E-Lَ��q`-�G!X�ը�F�k�2�_8���~F]��Tbܰ77UU8"�"S���bw�Y���@���˟v����?K��t�����q|�����WwuW���U��i��i/TI��3`<������̥<O	����Ҳ�C�Y�ц5	,v�����9}s��
��Z�W���2�q��촥(�{�2A�j\��5�a��ћ�1_u�y����гe�ڃ��è R��� �{l�R	�I1`sC���q�chTއj^=gkX*8@�z����s[L�Ʌ�� ��3LD�r�}o]�w�$�$�s=��rT�ދ'j��h,B�\�� ���ֺ������P�w�OI��7��o+��|4m�q��d��$/�����[1>C��㧺l 5�=U���9�~�snl���Pw�^�(y�v���:L��}
�j��%��fk<ed~)���h���0���	!�Ml&������˶T��1�|7��M�i�)Q3(�Y;�g� >��f;hq�F�1�d�j����X?�FnYϱF���J5�8�X�Jr�M���$J9�.�����ig�����P�w��ܧ��'o<��4�04�n�	��4���l�n�Ҋ�l�Fl�y�z�K��@{����%RQ���Ŝ�.X��_TA����$������C�+t8�75G@U%��[ϟ��],��#���p?���]Dś0����ؤ塃��[Y����ZXS;��%�F.1E�ش�<7����cz<8�׫���c�Ǭ��^u�'�ZJ��{p�?��z�l�gw����'>���Wk���H�
��#ݚ&$ەЖR�bS�[n7?����)Ȍ{W�Ʈ=!}��h�4�=�jN�($�>�hQ;:��qq��A��j�e�,_h�u��&��t.�ַ�W}Z���|�;� �Jd�H�N�o�g��� �j�b����|�(���T{ᙛV�4{q�C�?R���n	�Z �����v%N�3�S�t��ĕ���3�E��t��A��Ϗ��7uKJ%�Y.��!���h�t�Š L���PCݭx`�!k�xSJz�a,�N���+'=���ૌo�d��j���Il�Kg�Q�hiG}�W/������K���w��8��ۃ����p�Hoߦ��ɛ4�~��������M��
�r�s�7���C0p�T��}2��N�6�y��_�	� EUq��J�9z���ŠC�0r�~�A�Th��z���ե�9�u��I�9�?���Z��%/���E�Z��Pl�_2ߦ��<�7�qo��a�ͪl��x�M�ӣ�P���Bh�5�����T��I$6cLCĥ$J�z��f�w5�}+��S��p�~���b�S3gIw�ŝ/���;/+��2��R�y��B?"G�#_��y��MI���'pI(*�"�b��T�v����Ч�ơ;��a"n<���0�¥y�նرc�2�P#� 7����a��0��uZ<�x����	'�>���+��E���d4�{aIw�DK3H1�x�3jV�*�J�����N��y��=�
��n<]��cqf����ڻ����O=�I�{H�勵���ő.��SWě�/����e���K�%��{Ϋ�&;6�Z��n�x��t-*�Hsb|+�X-C��\$���w:�Ʃ>ǾZ�-���͟1~���D�a��5cN�!Ga+
���g��U��׫R��I��
$�Dً�@dl��z��%� 8+�C�p�c��R2�+k}I��p95S2&Ab5w48�}�^V�D��OAz[-%�9$g�@���/�\��gOp.PZ�J`�-�bV�@��~)��F�X�J���z��zJ��{'z_��mKS#Ʋ�!o���pm�RF�80G	 �
ڠ��_��9aۈ /�8ZЄ�E�z��H��ũȓ����&C`^#��L>"�N�I�|t���,幮�?�E��@�:F�:��a8p�$C�C#�+�e��{�z(|u��p,c H�cq�*u��&e	d�M��{�|�{[��y% ;	f���#�W���zǚ��	Ķ��80A���E_̑��̧�� ��)�P�ϣ n%4�ti]�:%	����)�H��sF�ME]t�1�QQY��h��d6G�����{�j8�g_�2���Wß���e��b�����'D�����@]����{�Od��Q�o8��PO�� 7P��&�DKH�0��[{��X�'��'߂ʾj-�B�7.y��L{�,�=�|�i�N��s���8F�E�ǥ�����wW����������]�^q��}�B%۵Wr]�̌W����..e]��\#�t�����#�&q)������/����~��~�ɐ;�c'�����W<d}�(�>	C|N�<�Z�rЂQ���e��R�O���3o�!/i����UXZ�
�{�����M��0�I�\��GQR?�\�]��J+�UO7ǣ��za���H6�G�^��O�k��B�Y���<��r5��Yv�&7�[��[q�p�7*��5�I�:�D��̈�t}H���Ax������7�ʒ���ܤM�=�;�A��8H�Q�9�z�kH�n��7ыJ�S1TupP,��x��(	Lr�=Z�9]��N���;#�y���h0Z�b23I�o�fll,��bc�J�k�5�W��P�`O *�u�<�ZheD�#!�{��D��s�(�����Ai�b�̄L����
���o��D��]������2�k0���m3��a�$����E;���tZ&`�X�4+���*21�n��ߜhZ��X��ducb�v4��pEY >��e '�+��I=,�;<� 0/��Y{Y���6l2Yt���b~���m�K���/�.R���aKc�{����M�Jil�l��_z��7�zaU-�oV��D\�pA�l�c��O���~Lú��F��AXU��(fF�7��q�� �	a�hZ��� ^���O�KI�r��ם1�C��GV�|N:t��{����r������@�;l�� >5��3?�j#�t��͝yE�:4�c>��Zmj��̠���Ԅo�	E�(�Ǜ�W��(�tW8�A3c1��\Zi�t��^trl�L>~c��:ڃ`��0��N�����pJ�?|S�SE�J�iy��W0{�,�U��ohW:��z�����s�t���]���u\u�m.��Q�ab�ʎ�I3�jXMT�NY��S�ȏ�#������>7x[Z�����F�X��F�^ h�S��;j=��K�<ٙҷBn6T�p�,X�`��	�þ/a����X�ɝ�����n%&�Q�y6��sxy*غ�q�ȟ/豨̙v����~ώ��7e���4��D6 �Բ�\jH�)�<�`�q	�Q-�fn�����t�P	j��x���b�dr�\�T��g�vx���£���^�sp�	y7l���ǋ���Q�n\�)ʏ�Qu�]s���Y_���~޼�մUY��Y�������Oۡ!o�C����Pc駫4�p��f�['�9�Eo���}n6�G|]v@�[���b9Jg�;�5�\d%N�a3��V�TM��Z��� ���e~�|�ɮ��2����;�㓑_mA�wpzbY�p��f�]��J�+�u@��'#�� �nF���v����n�(�s_5�+9Qw7@C�B.�R� V������EmB�9�Ϊ�c��Ӑ��u�� ��"쓓�vg/
h�m�o�H�������(�6	�	���W�S�9~�PdTlm$�o����b�������[U�,]��Xc�[lK��y��T���m��40�(�n���Xufeې���S&3���}}޺���:=8(��8h��@պx�yV�S�����H|<J���5诽g�@ wu!��ɡK�!�d8�/7�u�|�N����Bӗ\�~�e�}��1����g'���@��j&����./?�Y�G��!��gst��E��W,'�����pr�����G;��,D֧���%�w��Y�K5�e5I1g���*�)�Q�_$�$F@�
��[2&������������n[!��W#���&�N�Ӯ��2]�=
ul4[
�d��︰>�z1r�X�Cv`�y�UA��X�����V��^�:5/\qg0���PW�`V�MhK�J̆�8ҘX����z�3Z�"��dW�R�FdL���%�m�%-�o����E��7W ;R��OMFu��-CÒ��ϸ�m�AJ�G��7��bM���lIrf������(;�A���J�K#B)l��5��7SP���/m��$���� O�@Xi�Eg�^Mp�$��ɂ���������|��![�,G@��p����h��_Ҙ;}�`?�o�P�/iL�����n]���Zg��/ز5���U0:����F�I�rh�)���)XC!!��͸&���<�mw�oY��=_�?��)4h�'�8HoC�
ų�� �_,�� Y�g`��|7���X�Hc��Z������G:�����c�X���<p�	�F�����Oi  ���`�J��7��3{>c����f#"ŭ�}�s���R��Ӧ��ۇv4X�~�×�<&��Y�p0��d��g�!fɅ`��N��|�O�_�-�q�z�-�2����,:$�OK7$��u���Te�r���O8� c���w#���E������=Q4�~���c�Rݙ�u�	L��=h� Lx-�2XY�.��ݳ_�?�6o9�A�s����z��<�w�z�}��z̽W�%|%l^��C�ZE4�<��Z�8d~�q�_t�����/⛎?�0�c���?nb�W5�e�p���a��x$�e����������C�"4��l�"x~��#"��H��/o�R��-3��x�j$G���{p{�@Ve>�L�M��kI�Ec�F� �����?����i�-7�+�Ҙ��1g��yl��l���a �� ���eI��9�=��+�^1�h3�E��jG! w���B-/QEoT����隉j\C����Q�(E����O.��s���ͦ��N������(��ݍR~
�P�����ɭ� /z���MPO����x���R��1�w�G|�s��#��_wnU��",��]�Ng5Z��F����55�HG�j	X�����iA��p/��n_��$�&�6�����%������$�;�q�.D�v�Y+�Z��I[,K!y@�Ǝ
�%�lؖy��b��4|�N�c�{�4Y^�˪���oQA��%t��`a����*}٣-_��x�׽�����S,{��}j}E��"�4bk��4J,@�Pg����p\���:�ո�@�1K��Ss��m�q�
�Wnh@h\+ �c`P�Y����S*������L<h�Q ��՞�N3����v�I����ms���0�%����T)�E/^��*)GE�t�Ì���g�mT3#�0�3�&,\��dFg�&�����hVB{ml��m�g��6�~�A�̯5�j��f�P>6�j>���׌�F���<�A��F�P�Mr��M�q~�t0;HQ�-����.c9a�82P8�A�}�����)iV�`�bJ{�y�Xn�Ҥ��X���|��}�����o�+t�;��7��'��7�so������S�V��4i��r����27#:����Yl��g�3���~j�h�"�CU~�?�>���������S]c!�����{:�>��^[E��x��Hd��|`R K8�܎8�H|}����m���u��rG��ם'�Q�e�lLD�x�?�;�}���Bk�{gPN�����>(aj8� �5�?�M������� �G�NL������ɨ����9�D�cޙ	J�6\⋋�NT�B7����>�2���{�����InӬ�����zb5/,�f�{p����Y۩�V��ӣ�J����*��gXz1z ��R����{Vg����<���	��� ao������`�&.��:��������M���͔n��l��a@���_.�)�B���~�uy�^�k!�x�$i�y�G�����!�gF�m�~�#�E�(L�d E��f&�c]����S��|V�Pw�}����	IQ6�,�v�}���
ĳ`�K_����<C%���o��4�+fsV�v��f�Z�78"�ʀ�a��5w<Gy�E m��p��� +�	F���촉�$��D�� 5 ��U�Q�Jf ��g*$ȧ5��y�&$�P�ɮ�4�wۍK6W��:���q�@�ߐ����)]�w��z��@?��%k��pB>-����Ly�^(��f%����^�}����K7�����Q�Cԡ���ӟ�Ű4�����U��ע�	˭0%����d7�����~R��" �j�Z���0"6,�M}o�>gxɣ=}[RzZ,��m����v�c�O+�{���qAgwͮ�2����I�Q�ƛ�"��"���1���5Fw�jm������x�v9����"S��Xʫ����^ґ���j.;�L�/�]�Y��j盵��Q6��Ҝ�W��8f�~����E9�on�F�NSo'ɋ�
B�(Ӄi珗�/}g��;�eG	'���f��z<�H3�k��h�rH�����)���q��pI ��rSmh�@�(���1ݴ��.� X?�¨,�L��}Z�d97�hv��n8�E���D����R��^����Mg�I&��(�l,��䢞IkY K�T����IIhw�2RZ
��1�.�I��W�n��bX7t��c���P��߲:�V�U��(���e���X|�?3l�$Y�~�a��XS:���Y��20��#��K��O�:���p=k�����@BYb�`��n�f���8FxV �fZ�ʂ_|��7��@�27Ƥ)"���hO2�(a��S�՛��pg#=p<��d��b�'�I+�kы׽h+�r�*����0(��9�6��6B��?^��GD�P��%զ���k��ٿ�RC)	~�>���s F$P[YCWsʬ�I��9���t/2��њ��zV�c:9�mVZ�t)ɤī6a�W@a�%>kΓG&�
�L~�)�!ڕ0D�t�)g��u?�ݑ���Yd{eM[cЪΑ��J�z(��k/2����cڪW7��p�l�P��Ԋ>J6��>���$�ӧ�^j���
�>!-�m
f����i΍z���F�٨!V��Pf�
抋����>�p�>����?y̿���Q�nY����~���4�����,�g�I>���i�bQ�Q���k-\��g�rCx�;�/�⟏f#]9��p�,u��l衲�>��0�1%O(�<4(����dܴ��ݬ@�*��7eT��פ`��`���-���L�-+ݖD[���o�Gt�iy��K�JS��Yp�T��Ǜ�"��C�)f�-y͗\�G'�g�<��q��������O_�[~J�7~w�-�����lU�#���X*�Z�����N�""�1U�՞ی��� ��u�>�8���)�38_��ַ��` ��z�� ��
\t�_����`3E�g�y0Es�N�;�&kw#"�Z�z֓�R�E�3�i��$��g
�<�s��7���-�qG�+Q%gZ� &A�4�Q��<��:y)g�)�t��E%QA�j��8x���z^
+ᇒb�d���d��!P�g~f<��>� ����n�}�G�us��0@�����],���@\Z�`�E�\�p}o	u������a��z�����ֳ1=s���o�<��¥��M���[*%V��0t�W� T �p�x�1��w}�L��'��]�*G�b���T�F�h�b�;�)*IT�I�������rBxf��.6�>}H�L�/���\��_�}���<��m�/˟k�T���N��ż�
�����[@�\�Z`F�4[���q�*��9I���+��K	�]dS�z���"������6���{Α�V�)x*gH%��$s-lLܢ=���4$���)bu�a��OYg�y)x[����Y��_�j�gO��6'����y�>��}��c���z�X[�=��]Q�~43�r�Q]�14�Y��s��0�;,����^=�n���Z{�?���T�<���9.u��A�S
:wj�Wb�z��|e��?s��:��@���0�;Tr���ܛ�sjX4SsM���X�sY��o�D���4�gJz#�l>�߉�^����i�l���Cf��$�y!E�!?�A;�5Sһ�z���N;�W�ELZ���O�s�ǋ�%��hs}��}��<�<� ��>��@߶JM���!�D�]��~���k뼨�9ֳ,=}uB�X6,g��?��T��x����l�=����M��:Z�<;F\��w7m+�$��z�^�:�Ap%>$�hP-Q�C�H\!��k��I�=�4���Te��xF���P҉�jd��ly�@�ZuB�q3Ln2!s�)J��X�!0�,��yNw��a�g�;S@7en�m3�v�vl�Vqw���tF>�WX;Yg����j}͇
�`��Ի�II�.]}9w��
iݦ-{�AX����i�z��Ʉ&�h��nJ�2���cK����nw�ƛ_����Rq��ژޯ,�YQ�	�r�g� 9ք?j�B�4!p���xH=JX������ڵ$w�(a�k�ή��V�c��x�5� �Jeja"�oY��/X[]�����o�t���-}�G9�y�RDB�g����, _��ѩ� ���k����Cq=�͎Z {�ל�<���p�R�t=�:v�� Ԙ�9:�f�1T"~����[���V���slyϴ����B�O�TJ��'b^w)�4�Cw��� ��xN6�ˢ��gȋLn*o+�ӻv��LRޕ� �)=J�!�WF+���?��Ṅdv���-����eʛ"��5�A���B`c&Қ뾕��{�ʿMG_�q��.��k��+'6��c�0�S�r���+�� 5Ӏ�t�������c�4h�������ͷ��
����	��R=����pD֚h����U����%|8i�F$}����p��rNp��z:�q��z!� 7�6R�8mm�^+R3�ha��[v�ݼ�Ol%�K�o������{�饩�]נC`s��e5���W'#��E�+>{#8ˀB���y�Xb�-E,�~�o��_3�AC�i�eYx�ڿ��17���47\o(%�~�|�m��� t�<D��q�%B㞘kU?nO�34�ȿ��^���Pe�_��U'��}a��+�(���+gG��J XIo��d&�k�Pƃ�Qa���8`s_�� C��?h��{�\�l3�+��.w_�A�$a��(A��� ����{P΅`���}x�uNg�+-I��KO7��1��7Y���3�P}V��6�}�y�߰b!�#~q_���tE�FR���qQع�7,d�Kܡ}�GbE�9��t�"U$h�ƃ�pWWzU-��t-�� _k���64���X���U��V6�| g6�"0���<�z��Ц�w%��qU��HCp����`S05(�p�~M��=tS��C�n���$�5�KHeH;
���s���)��%b-���o1�HaP�*�ۥ��W̄� ֶ] �3�o1`Q|���- 'ο�<rpm��/���D���j�6��Ù�8zcx�0
����e3��IgtC@�S�!��؍���&���B���T��FȮ٫t��ϛ��>��h�������*r�xyzt0���U��:w�`Zjc�����@0�ܫݑ>ǂ�ѐ��cC�V���*T.�waLQ��ݎ�����5Tu�L*FY�!q��?��6r�ԥ.Z.����+M��ӟ���Cl�p�������j;��T��n҉&������Ӑ���3�%��q��c��Ő��z����_^ꥇ;�K,v��=���x77T���r��E�� �����&`yM��K�tC~ޫ>�����Qz"�XN|����˅h_�\�e���i��[����:�ǂ���r��H�د?-��[�ng�D�{��7���CܸP�kpgL���-�"�ef�l���UY��~�1��?�1�Qp�̖g1����6�~N眰1���^-��g���0�a*����j��Mi19�K�i �ҧ"���_�Jt%�*����0&��4aitg�@�_"���m���a��*��d��f,#�~[5�9DS=�!½pPH4�D����p����O��(���}��s����f�Q��}	���g�Y�ߧ�qc���j��:
F�X�¢|eUOw0�,3�\f��%^��HIV??D�ZSnjc���9�U��1��Z,�Zw���ʫ0���~�1�t��yC��`?O�y���.Y�e�tߋ�����!�]�祪���]��5a]�"ٔ���j�wOiy,@�E?>< �8v(���<=3��6-��u����J�Ќ�|��NA������ɉ�`�jG�W	:�p0��i�
�T մ���V��E�Z> ��}a�G��D����$ؕ��5����ώ0���16��f����/�緼7NAO��m�=��}̗����{bǆ�[�� �~��)
yc���ߡ��O
�R�}�u�^[�������t+2��K�R�i�A�657�20���Ji��nij�eu�v�
�M��SM')v^����Ղ��섽����������o�s���X 4������s�������j���O�Guv-$;�{|[u2��ΰ�����rV<����`d��齵Ζ��-ѽ�������@3��U�5�[��r �j��^���z.����*I�|��A)U/K&l7��/��{�������lGŽ��n��39f��	A>%{$k�?��j~M{�O����Ke���Bk�N�Y��j(}�X��R �YVM�CH]������E ��쬯�m�o`m����YۑMEg�Cp�g^���|w`$U�H��]Oc������m�������O����E��q���{$�.���b�@s��|;�HE���P�q�B.�<�g��,x���uG���q��!���"��ļ� ������E���t�U�ct�ʙ,��̞p����_8�>}����	M܆.��v���N
6�'�M���$���&"�E�>�8��N؎IJ�?A.���)-65�5E�8�4�ߠ54OR6�$���(�w~���%��IHc����d��4�?70F��2�_Rϲ��Ƚ���$% ��o��^�U_m ��𷮐�J��@��� �����~@~�?�bI�h�gY�BI{��P�_0�
��S*�f�]ݣїfO�Tfw��|4뫺��?alW�PP�cch�����C��X��@c��^��P~����K.��%;�V,�Ȋ�d�9~E�	�#p���)��з�?f|T������Ҕ�9�ҳ;��ʿ&����o�T�6����{�걚"Y_�*'?��ya0J�w��3� c��uq:>1h��yE.�:���o����b�t�{�{�=�Ɍ$�,���.�,������X�tZ��'�'ݺ?k�aB)����![�8kL�yx�z�H�,ʕ�z�e��l�	t>�2wR ФwV<B,�`�;��� ������=-mn��*ڧ�s2H�}�c���9�l'����O4c;Q���fy�:��iԧ|�q��4��jw�>D�O���͖"gţ��p�R��3��s���2N9uۙ�9��DAK�����dg�=�|��+-��f�YhOX�O]ϓJ\-���/-��l� ��Δ1�s���]�]I1T���,֩Cy�"͘ج׌�|r
�{!�Mu҃K�9�A�u@��XI��I��_�į�,�k}8[���5���W�0.�^I��E��~@Bػǡ?�?_�3c����F�p��D�Ï
�#^�%t��:��>���hޱQ�Ca��
�'�Y�,K�l�"��1��0������ӽoӜd>���������uE�]���<���VO��Z���qS�B�јI��1�Z��:�p�j���E����RG���_�8���W�H�ȉ:�[.ł�QZ�:'�YB�H!d�7�l^L4����E��9sP��!���`_4ξ���oݞ�� [�Qکk6n����@y$P
����p�cM'|!���"}͉^�oxm��-�c�ڼ��r0�()r'Lw�!^��ՐcU�5�|��sWC�}�*_-I�8��C�#^��/���»����(���viJ�����!�,%�������_�:���_��ا�oT}�|�/\'j��ʪx�N�K�u�!��5���Z���oF��i��UI`L���y>r'�ĺ���n�)��e~ȕfr��S�9��(s��RF���i�yGd4C��f��Bb��U����v0xg�T֘>��kK��@ةa;�9��(�}��&�R�Hs�;�?�A���+g�2b�V3��a���$�*�5 dX)��W�?��O�7`�M�ֳ`�+CI�uB��/���}�ݱ��������_�LϾ�%E�[5�G�ٵ���q}3U�WpR*��7 |��y�Vƞ�WF���@�
�Z2a��5�\�HW������Of����ͤ�;�#0����t$ 6��пo��a���+%^��,G�ibQ��+�7��,��ĉ�d�`���|��:�x;qī�茫�Y��W������71V��o�<5�|��I<���D\ ������=i���*r2S�!�I
�aG+y$D����W���(kXhjp_�!]X�Vk ��T�B�W�h��J沯�:�^]�����d�|�:s��V�T��A�\q�s�T��Kѝ�;kM �<����ߕ�"e�3
g�p`c|2������
���p5bgu[������Hd���9�lt�e:��J ��s>��q��}�ۚ�2D�����N��]T&U(gv����3�����ŧ&=Xl����8��Gl�	�x ク&�A��RA���?�ʅ�p�лC�`��@��c&\�������^Q[LS�(Q�=���2�g7ƲYiWE#�(�tbE����ۃ�e�|	��!@���~M���s�鹬���cq�����5��Nكۣ?����<�;��?��D{�Wd�Dx�p�I�̡�����$�;�u����cRb�����ŻHmKm<��1���$tz�\.�,��kw4�:������_G�7�-���+�vC�Z_�z̷�7��Ͼ.v�q=hh�tk��|Z���_�G��t%ۄv=�����LNƸ�6pf#��?����.}����P�2$_E$G��$������=jŋ��]R
^�}پ�:V�R����?8��\y���S�i��#�z���W�C�syis�����g���N�s&����&	����˱�ʭ����1�����x7<X?ݕ��glTǣ�'�.O0�	�
_���L�?!�E�i��G��|�I aN	X�B$�}̪7g�]Ч.�50	ϩ2��d���ע�ꑎ�cF��*1�ʟ��`z��m'�L:g�jj��7W��zs�c�OdJe�ĳ��gLt���ϙ*V�
�'<+�˸3&Ҝ�F�G{��^	B���_�D��|�9m�ƍcM�X���m'E_<H�]I9B��,�@�����Um�d�'h�̒�;I��)$%\����á$�b\��m��b��%��? �>��>� �D�q�{���EpB��S@%�.��'H�'G�S��ҕ}�1��KBP��}p��h�R#&��KN����T	��F��=�L� 58���ˁ�1�5�o�T�N�K�e��b������r����L�~�N��8��Ň�u���+��V+��� �U9|(�_�'Y��v4�JIc>�4�0H3�,v*�m��cA�I� -�6���E3�u�������Wi/������m͋H;���Z�C!��d�Ű����e���O��e�(��7==Lx[) j��^vT/��@���{x[zC)�~u�5:���PX+�D�ϩJ�j�N�xu��n�$��͵�ȱUy'[���\q��ps����C���'�����O�?ڨ�k�[�,/E�ϟ�>~'�7����-#+E ���Ǵ��_<��iUm���{;���0�\�X�*SU}e(�����Ֆ�{���v�Xv �WCe寥���:2�ԍQM�B>�i��b�L��&(�l����]����0獴���iP�wD5N{�Be���I�ޔ^�ue}�-K	,����}.[�sEd�a!�� >�Z���W�
�>n�����Aj�1�қO�|�e���Џs۔/�e��A���x6,�+aC���\9\�/E��ݞ������Z��\8���)`�o:�=8��U�\0�lȪ���9?�����h�J26��H9����e'wV���EPm�9ƘCD���/��,V�N�[�kď�������߾��)p��i7��!w�ת2o�hf��NQ9SG(>�"�� ^
���mɿ2��<p2� N���3� ��g`��~1T�1��ajSd�%��dG���$P!� �x���\�1�3��K��[ע?�@�7l�m�3���?�����}#xd�~^�	5g�g��P��!	�D�e6�TE�xn���c��0�xCi]����WS���[}�|�����y�+�d�D���F����
��(h�O�9v�*�C����xe��p,'Y�i�T	�U���V�d�=?�G��z����^��!'k�Ti8�f��!�H��@���k^����C��貌�M�kh�P��������BD�#$U�^r��#��w�$�k�z{�M��+N��<Fp�)����ɰ�^0Bx�w�J�cGŻ�	M��~hȇ��~�Y�enN�.��F���cQ9r������[�ys9�țin����_5�ciT�bgwk�Jw�C���j�G��6}��sd�7n�9?�Z��!B�k�*�m�W��V5��/�:��I��T�0��6�O�����.DY�T\���CWm�j'(���ߟ������-�����u�,$瘾�u�I▞ף���Iq��q�����@1�=>T�5;���"�~��}���H���ܽlU�w�öp��'���V���2�6N��]����1���V�^��C�w	Op�M%��M7a��d��>����S�$M`)_Lra��`I�cY���(ORe;�7%��6s���$�P�̓�:fN���x��?�c~��E�v� c�X�-J<���lU��q���\ c
���d��6��Ô�%�M�>)w�ox�����u�;�h��PD��l�>[m*����������W��R�����	u�տ*�(��T(MBe�$�2���`q[�K<n#�Ŕxχ{tp���U �)z�7�%l$��R�����}�>7r5,,�#��vS��D����w��0�����C�pKϺTK��	�uKyܧg��A *��(���]��O�u�3��L������ݟ�u��=�Wv|l�/�/� Pfws�����f0:6,@Y '�JÎ7�G}�UDЊY-~��2��;���(�D�T4����:��@AE�ӯ�y*��"������g�!/�O��5��N�U��)0��G�ɖuj�u��Ǟ���g4;�j�'E���n=�ب���-3�e�O`����nS#�bƨ%SF }�hsi��}��
���"6f�6U�4�gm��g��;I!|ّ�JI�z@�����I��(��b4VeYoK8�z1�M}>r�_��TW+y�a�wn�O�n���&�za�J�^@Wƭ,��e=�8$��u�T*�����I�c#�CҜh����ى���|���~�'��p*x�~�ˑ'�"�&����߬H�6_O����=�]$k�N�>�����meV�(L��L��l�t�ѥD�<2�rd�G�<��\���h�b�xЈ	z�vJ���Yzk9��h)W��q��j��L����͓r41	Rac�6Z$���X5�8����̵]F���?���Mᇙ w�*5[**��e��E�����n˲�gT�6eJ�#�{z4�^�UG��T���v2�7dbi+9N�ӏ��� �H�;D�&2��q,7Ҹ���4�%��L�?ʀ�8f!UY�hɕ��{aD�}Pں_�����Y�d/���>^�a��{�w�m�A��E���^�b�
�����΄��2(Q��@��$��~?*�H-���-�=�d�Bl^#�?60����"�b�?�Y@Ε�� �|i��V��V,ǳ'�p�/�ؑG��R�Z�;S��oV�:ڽ�O���]����è�ٮї�uWo{`������U6 0��NY'�~I��9��{M�FW��<�꙱ŻT��a9l8�8t�İ�����P�:vx��1��cyQ
�vd���#u�������HS�zG�V��ʷ5=�o�1�T�	�H�8��û	��n5Ѣ����Z�v���f���y�O����pIÇ�OF�S�?�\�ޚ�}$��^�P�q�n7ޔ���maOob1��W޶M���w��e�v}�GŅ�ԉMtȝ��y�*{/c�L�뽔�J�.a��`�r;У��'��15�g=��+������ζ����*��\���虥�[W�e<i!�	��|�v0R�����)�ðLU��Ǡi�������ө�[�@;�y�A�a�{ڝ��>R;�IY>��>-;���9�m)�=,�	*�o��:%�p�F�������I���6�����']vcz3�	�&��;�p�'n4�T���Z�>���%_Ԟ�@�t2'}T�Z$^uv.��p�;!	�"�4���]�o�#$�ӭ����D�u�]�c%�@��">�a������Xi���X���{Jr��B��X�r��p�c�kG�I���� ��]S�[峧A���[�(�PQ[�&�j�B�7+ ������2�D�YaU�;Xu�2���%lhS5`y��34ݍ7,���� ������z������W�z� %'c������}�
º��O��t���u��q]V��� 2_c�d���_>]+���x+N�����]�"�D��9G�+Y��/�� jֆ�`ց�E0S�"�ew?���^4�����f�b����n��UH�G]t�tμ����y��9���>ʊ/X�
�цr�i��RNt�:g1\W�%��c0�Fl)��MM*�`&"iB��-q��UN
����$w�M�~܌R�y�a�1w��`�&A�C�x�n��������3g�����o�{���e��[=�ux�t�a3�-)į�iĿf�P�;�����(�����#��q�C������-{]��y3�?�Z��V~������J8��>Z�f�;�p�my�w�P&�t���-砕�/oPN��w�wS@�x���v�|:��%*��ݰ��:JkG%��j�`�����*o���g�%[���<�n]_�w��+��a�*s����\���OY��α�c-��g�ev���z�}��r{&��S�Rt���bT;�W�����"?WO
d�F������>1e%�؇ �N�����cY����cŧ}ܞy�:�-�7|��f��Σ���hL]�o����`ʰ�d6/��L_qPBP��\�6(PBeۉ��3J<,��0R3��Y/�kO���Uy�)��$r]G#ƉD]	�[%�j���B�PL����N�'r���y3�騯���hL�8��`x(`T�ӝͼ�]�{ο�
4C�ɥހ� E}�I$�=�����0�VEDLdz��u���Eug ����P����؛�*f��*�b���1����fGh:�N.�`��x`��ҁ�gz$����b�RǞi
<��;M���y��}f��%�Q�~\(�N�ҥ�9��*�(#��v)�SZ�fR���(����c��� gCy��,Ug��6��� F�p+��˓�ƤНȮ��7�dZ���Ÿ�rIz-Բ�L��+6�&�� �~G\��2�"�D� 	��I��a�%L�,;RA^�J�3DI�_Rhr���eG+	-7�U٦g'ş���hݡ�`��Y?&�3%P��6l2u��b���<ޭW�!�,��g�*��|F�� ��|�w���Cn���sa���U+�҈��S���mB��+�g���1M	'�x�ך�������!c�}��>6��(iT׼̕����섾�F�ߡ�T�ʑE���-��s#�K& �*�EeMe;��4�uжN��[���-PO�K;g)B����W�?�"��b⍻�Z+�44�����̏�j�����ߖŹf����4�ͥ��鯧|����*��C�
�6c>oZ�b�"���nE����ٲ�{�����WW��Z�.8�E��M�˧�b�Z6���GS�Q���!�`+�>�!��.�����MYs4��d`��7.�x�D,~=�iu<�TR��evq���
�k��b����L!��[_	����AZ�զ��w<�X�y���0`s�B�Sb�ӯ�b7��}�	�`ϤȌ�Qt�qM~m^��V@�d 9�1BH���)����$��(5z�"�"R��hQ:DJ�������9羯�|�s�Z�㒮_�S��md=YC�WlӅ|wݵ��y��*J����4B�|�&M�L�&�U�~��mj�k�j���ږQ�����k�&Nt5�Pz�`��+Tѩ<��$��qOc��O�?gV�bD��^.dRr��FLlT������6E��|y>q��hn6�<U_�u��{��5$���{���WHGk5�,�gWFV�10��'�1�4�K�Iu��XRV������O1/�)9�e����K)vQ��cs�I"�X����~S���U-���r%2�Y�����Oͭ�pګ-��;��������� &�[�zR���/�T��:Ȃ�Z&<�Q�O��6��?S=�*�C��]O�-��*.���DKF����7���& ?$��8x��C�@=^Ј�$�����?-[v�N��"��$1-,�\�[G}ϖ����G��G�m�u��?[%��o���Oqe��$��Jh�u�0o%�۾<i��՛��k�kϴ�q+�����D6z�!�)h7<u�/��������
�9�FG����)q�w�Y�������g�ζ�3�ӗ���Mf��)����bA�z�����R�#��Ѱ���o��ѝ�*A��"T[�<lgZds���h�[:hkV��PJ�+�4���~7͞xQ�-Y��ю��vk���H%y�:��L+�)�Q�m�ًl��*�������9s�/�7������< d��}��<�DT��!*fPs�vd���I�l
E�Ҕ=]B��x�O2�Jz Ŋ��z�q��$xkI�ǻ/�iO�/���ؕ��}"�0M(�%�  �����Q�5O��Hk�Q�~8-���ڞ�&RY��%�C�k5���s��Ν�������?&'W��B<�bT��[�N&	�u|El��q��kVK�u����bV���%m�K�X�)�ƽW1��}�1ĚDq���Y�U�nN0!'\�	Ǽ�ѧ�E�I�Uu��O��I��H�pfӊ`-�C�`����|߰��ʚ���ߩ���������*�V�`1e������ֽ�r�t�	t1<�n�H#x�+�ǟ$?1K�ʄ$�uՐ6���.� �`�f�t���oy�� S�}�i������M�F��,�Wup�q��Z����� $r��G>?�\BjM�M9�R�>�V#P|�[���н!X�m�&|WS��L`L��k_�p	���N+�| �|L���J��u�դ����n�0�`~,��(�3�����)ɭ���fb%T�w皆q��2im��_-�<�� k������mg�Ly�Ⳬ.=����"��?�Cvv�����hA4<����]co���w�0�38�(�iq1��U�Gg����2��rs��͗F��q�T�������5��3k����W����� }��H�٩ՙ*�]AY�jU����r�ðy�$�eP/;�!�=�*�\w��ޣ�+�"��$0���;�r8�6X��,�v#��~�!㜺����2
�������S�<���\X{�|p�v�E<�	�U����0H�z�T�/�4ݻ��b�y���q��폋_o������,�{:�9m7�h�o|5�2Q���m.<��q���>�RO�a�f��y�_�Nx���idPj�^�~Xٱ�eb|_>xA�Tߎ��ɮ��?�D$��Y��^( L�#XI��o`�n�)=��%���U4��O[�����7�F�XM��m֊����S���y��Ig�7���zt�1��i]|Ⱥ�eu10���ÕM�h�t����Y
������C�>Z>0�F�?l��-b^�&k�%�n���!+J�B.�����q1�o�G����Ucx}{_�9�f�"�b�rչ6M��`�$`�Ʈ��RdM��S b���"�}�.	C�(�T��^�r߾�P�'ZRX7�^�:��}gO��K{����2@�K�:��-����~Щ@���f#X�t	�����`T��MR��$�SD���_��D �t��6_ ��{*� ���܄t&���̎��y��p�&����U��x��+.^~@��A��雟\���2( -��p���k���hQ��z�j$�^C9���+�Sj"ױk�W�
��hk�.�s���1�zS1��U�z��O0蒂ȝ;d�6�T�YC2���L�ҿa_��3?4V�^I�!��$����S&h���B/l�!g��bs�P$G�4��5L����.�
 �j2�&��{O.�G�=�ܺZ�i�5�kF�^�7Oh���z��q4���ʋ���i�y<�t��([u��~�#ڥ�H|ĸ�s�!ژ�D<��Ђ�*�����4}B�aN�?+p)��=s';�F>�
T�;�Z>���oᒞFk��;��y3���;Q��F̏m�Ǔ�����)7#*k�D��h�vޚ[
_p��5��Ͷ���pd=SLp�R�"�c���-Zeį:�(~W�{� ��X�<ԁ�m�	_�q��H��[L�N9�HzhL��.�1���~zЧ�X�	Y��!��]1�<AL�ݸ���.:Ka�X\Rr9�I�+��ǕVnqG�`m;��b�/��#d#�����ގ0$�^��y$�b �I{�h�3�/W󽀉�>��HO��iۿ�i�	���<Ԟ/.�^;\k+z�2'���{�?�oD܍tQ9��$3a9EGJ`"?��~�沞�F�xP��>��/�Ei��gQ��w��9����~Z���@{�C,
���ƣn܋�Dt�m�i\+��! �X��"���b�"�M8��G���ʭ/ɢ��ٲ�.�t����|R'k�a�̒�~;Q,(u��_���R,�r5��yy<������{B��i�3��Sf�k�-:ʿ�s�y�n�'�h��J .ouL��8��j�G%�`�q����,,<�ޭ���.=�����zvr�ń�Hȇ���{j�aG* q�p��?q#�O�*4�+�ՆOx7D���aj��E;��ՂF�g�S�eO�42�7��
t%���i`��Q����9���[�	\��N�мW�ɔ51�Bo�W���`��/5�Sjc�g�G�#G�7���9s4f;����5C�0�s���D�b�v8N�{�F�7�5F*���k����N�a�.���J��},.�l�w5��X�|��w��{|ѥ9K��8���Y�C�|�60	ݹ��g���,3<|K��[��t�#- R����o�3+�$�Q�Ռ9���3mT��%��*��<���s��nf�-�ׁ��;x�нJ3O>�u�hgn�/K�;�wz����DM�"�P��a��c�i�Wd�,�s(L�-�o1$��qF��Cy{���T���*���?�rP�.nƣ�p���W�b����0������^�8KK� g���b�N���K�Ti>1� �=�bƦ�Xsm}����.�nT�{��
Dp�By6T����:�4h ��G�ZEuD�FxJ�'*�T	6��������{E�kח1H��z�.j��p��]�u�S�����_G�ƹ�O��
P�� �d�0���f�I�A}���vJ�>��$��|1"���\_z�XL,�\�1z��ƨ]�o����"�^�P]��4U���4X(������j,Ƶ��r�<VWA�����R�?5�V�v��(��X�'D�zx8H�  �r��J6
$L��*�[k`}��4��(K)k�a_ixJ����Ҹ�"��� `]��TVRV���mv|�28��bY*a�_�h�@�E�z7��%<�ѡ�.�G�2O��+�S�ۼ�庘�M�0m6�d ��1T����	��f��i��EXg?�^li����̊@_?[|䭚ּ��v�}8�Լl�� �ED���f��_Y�L�������
d�yy��?%��
5�W�8��k8�?��V���AS�v���k<��<�Ax��T��ʫ��� ��D�v��[^.&^a�r�j+y���_ؖy������|��/g;B�aԑ�Q��9�������_ij��T������u-����M��������ڟ�ѓ���1/ w+O0?4�2r��l�|Ѯ/$�_��L���H�j���_��Ӓ�Nߥ��-v�;�39{�Zˣ�a�=b$��W�P�0���;��A��Y�W��q�&{��=,'���6�^����sޙ�=�0�ۏG���{�2ԺmI�����|�,�d���z �:�cr����	~q�H��tĚ�/;?WI�?@S�&b@��l�X�왝,Vd&���}yQ�3�����u��5���X_�I�� >�cj�2>�@w&C4���.䒪�3����Ţ���i�U��M�/`���٦_�_�>�����_��ǫ�7��T���;�Z������wS��f�瓶��32����,�`�GL'���%�^����l�kI��o-��۔�7biEL>]��Z1eԣ.Z{c"�v��z)�!�p���b��{�A���N��Aq������hZ���Ǜ?���t��K��
p
����5aW���Y5�@� ���%����a��p�*�ᔟ�(�^�>Xar��Cs��Xi���t���}��M�d�+I��d;cݘ�vr@YGj�=��u���B��e�ġt�C��mY�c�P���*qG�K�e�ף:��FsW��zm^2��zq�ď���r������~�>2��9�;��v<�;���'�l������-�H�l~�1��0@����E�"��HBlb(3�_Sɭ�s���4������o�k��
�
�oud-[�Wُ��h���NQr�<��y��m�,�ʂ����ɤ`>���l��I���o_ONF���DY��h���7#�gs�?��re}&���'F�=Ͱ�\w�<�vm�|�ԝC�si�c�ZXtߺo�m���+o�c@��`���P@�~	����+��Ҕ'5�Yh��z���[O���;��G��\���6i�������/Y��������Rrc.N��<�t�x���ğ���s^d�V������+��#�G.kS+�a��1�%?��fd��NHk�1�P�e^�ڟ���sW�ܩI��������ߢ��5�:���I��J,S�C#�BWwv�L��Kxz8�J���h�0���_���'h���S�ѓ��2+]
���;H}W95Z�]2�|P�[~g����DEB��^���;��_��Pi����|h꒼�|f�����㵧 ��k��zb..��?(�8�dB�YLen��s��|}~=P뻷���=���
�,��X��1��~�bm)�o��:H�^PN���RN��;N�<'I���Z(�*�sM���P�I��Y����b���ׇ@	�`�%��uy����^`<����ú�fd��5�%x�v��g7��EG̸�H����w&-��@��2Xl���/s����[�ד	��P�>�ź�2�;̮,[<�G�U��A,gi�%�|�~7��9�ʟ���������+�gt�J&���U<�FHzU/�`���!Ų�Y��N7�)�n��4�ͳ+�^5ŎW~��.(�E�}��<�s�%O�_z�]:2$��× �k[����3S��^��|V ����/_�TGD���s'}�������n��M -��k��,KN���ݭ}VCd�C�@ [1ޚ�}�nQ�R��S�?����f�.����76iOF��ι?Y-���=�cm�m�Rb~3�>)_�y������K�]�M����
"oP;���,1��߅ӫ�a�}@%<�1�SP���F�������nкUs�rM��,�&5�(lZYnz���>��5�Z楞p����< �u��ֽu0��A����4f�R��<�>o@��
�Da�{�Ŕ=R�x�9���ɟؓ#D8�e(��^g�8H+�&��+d7�6u�Ȋu	O1���Ҋ��S�����8�[������/���D���T������߾ $vF_>V��Gl���FZ�K��he�WdIbڍ���ܐ4íP$�:�������h�JSg`�<՛���*��;�.
��ӟfD�=Z�����|���/z7s���C��I7�Z�XA.��k�ֈ�Do��̘���<.�=��.Y@*��Q�ӧ�N�.�oDnZcVu4�ti�k0���θ�s��H��}��u9��v�rb� �j�MTa����Ƃ�b��-�cY����Z7a���I�⎺����(@9�q&	**ݣ��]����'X?ʜ�q�d��E��(��Xt����y�m���z��1�:��m���,[J���V�>��沈(@
؈���W�;�����ϗ��E��KK�E�6���J$�s
K��b|�kh����ݱ@�����u臀9O��6ȿJV��>$%��zj�w�5m�1Zu)��LD�����Fw��嬰�u��R��O��(�Υ*kgר�@�FP�#��i���J��$���~��jE�鳎�+�n2P�s��Q ��ۜ�����/E�ߟu�y�މ���d�V ��Ӥ��1xft�E�S���/,}�/@{�*���=7P&;^TFӾ�,!�^p�2��|e��v�Stg�)d�K�5�Y���Q]�,u�d�:c1K���ʊ{v=}�H��e%[Ϸ9Jw�`}n�yf�"i�"���&�����9;$<9�j'(��M��x, ��Oj��=ݟx-�w���|����X�D��R��7tkE�+��[DNlJ_n/FH%��GLQ`#hl6�l��r�2�������$�M^ @v^���
ci�n�N�Z�C�B ؤ!��@��m*�-䶹�PN-�i�Jű�}���E�w#~���ör�s�vy�1�<�}�����P��1 ��-��|�_��\	�3���>�6t=�`�8� `4�[��`$�6#e�_vpw��Y�K�E�t�����������fHI� R��bP���j��,g�Z�j�W ��f�$W:2��H�k�Ӟ�tk��jp���aw��s�cT�'� ��Щ��t�x�6ќ�?Nfd��P7xg�Cő�Kװ�2��@	�-�?��� (]���cԋ�S�]��������M���3db~l\xʇ��}j���8@�k�<��P��x��L3��q���b�����%���͏��`�I�G�cl�q�8=���5Y�Z%�+�*�p�?i=�S���ߓ�Ez�Ƙ���s����K����6�'̵L�ݛ_z��F�-���$��QH�Л�ʒe�?�kȈ��	R�4��~+���Ɵ�/Ό�fC�L�����7�T7�<�?zl���|���Rv��a֕,E��k�0��#k�\-l^�V�����L�j݆�ñ����?���Smj)��t��em�jx�+*<�D�~X�>+��嫔*�����B��}�+7}.;�<,�'���Ɋ���؎{�7�Oa1�v@�����X������ʯGj'����i��Ԗ+�ق;��y9z#�锇��7d���m���y���b��Az���4�����&��1.KsX9���p��r{ƶ-fz9��쯶�α�T}���,�	�4u��Q}������'�	�]��qf�~��?��s3��E�ƴ���qqSvLƁ�1��?<�I��cv�b�� ��(��]RD|')3�0Ѡ� 4�gZ���{��3����t��JnLRm+��{e+ň!�\�F�䤁�0���y~�jWl�f���a�O�E	˴����g>����V+-'�/a��L�)"p�"Z���xz�ބ�q�_�ǫ T%�Ѥ-u,��m����B��s��{�+Ʒ\<6ڿ�� ���4��Jf<u@�!����`��9��t+��8K�.�FV���Qo�G�N��u���8�ێ`XCT1��+�31PH2؍��dL��.ؓ�n��&��(���33,H�!�Da!2�֭�GV���U�����{�飔+�{5�~���v��)�L�4��-�6-��L^B�ؔ���ݺt0#}gq\���� ����Q�0ae>R_6<�h ӆ�U��}�|�4X�����R���n�f�K&�����է�sn�Vw�ҫ�z������qA�y?���8�W@�67`)ჽt$��ո3�)'��$}K�]ȏsrмy7zi�"w���6���)�m��� ]��j��p�i3�?]��]s�<D�j/�bA��%:~�����ė�����"ى���M;�&3M���h�->R�<`�>�hߩ��c�VͲ}�d3͡X�1���D�{��Y}C�8KMx�G�q�����4�w*i��R����7%�S����3��-,��sp�ɷwq���hnچ�{ڗl�&�`��~�f�g���[�ХI �[��/fL�:�DL��T���ֻ)���3�k�f��2�o}�0?(���ʱY�56��ʡ�{*Gᔖ���T��BRx�`��?M�׾	��]T���8Ei��E�Ā*f�):B�V_��E��6���ӛh����+o9W���/�}�/��'��DLyeq���Ԙ (Jai���6�m��x`���(Ui��qf\rz$�G^��8b>$� �[�D1
�U);*�I(��U<�1������ٟ\�N"�Sҥ�Wq7��p�h�r����4a{,���D~G*�~+�o$EM���s���AJ�s�Te�}����i;ʼ�|�T�wѯ�1T�O�6j����R����T�Ҿ���05��.ŉ�Ǆ,m�
�}G,��|�;��0DoMo��~� .d{4���-5�@{G!AWHF�E�C��\�:mc�&�T@0"c�Kp�O�sLDPA���_Q	�:.غ�aG/џ,�D�wN�<��&��2{���A& +P��X�*ws! V���R�2�;��:���4W�׏�%�,���$l�L��jA���/�Cӝ���c5�B�I�]7#��D.��h��p�q����g�r�VwMc`J���������n	]8_,��ϑ��fy7��Q��X��U:~M��	N��Wl���?ˑ��t�� �n[m�Y�JF�a#�a_o�H~|��l�a�\ 6i.��Ç��ft1x��6�^\�̪�2g1���d��(ln̅���6����b����>q6�t�ޥE��V-��,��xd�S>r6�	#����/���P�mM�9�D�Xl����� 
����[�����d�<s����|�| Ȭ'�v9��[7�a�U�>}I��zh�1Qŧ�?2�8��X�w�6�u-z{���Y�[�0N^8��J��:&޺h����yA�{��G��*�*��/�]s?i� ��m9�e	>6oմ5�����IvN�6M��f�k� Ʃ�{��c��+Pi"?��T�� �R��:�	�~�&R�.�#�X�������?��b�_WGҵxG����'Y��!�.���؛de��\��$�я�p��Ex�HOG�o�1�@c�D�=���EvIq���2��+�"a�d 7*Ց���Fg�洧��лfG�k�jc&�ͅ���E�V�G�]�v���T#T����p,(7��`�X]L���bֺ5���!�ٮ�o�Ƣ�I��{�p���������tv~�Ě,��9��.�6%�k�?��� �X���]$���ﭗ>Bo?��G��e����/��Y����R��K� t<�f��x���V���(*$���9����-ےQ7ڕ��M�@��kf�V��@�l6�yz
�C�f��R�|���f!�-?��	��
���r�}?�t�d�<R���u���MX*[��ћ�#��\/�UII�R��+�.L�la�h�g�������yw�&��Q8�$;��8�s'�Sp��Q��h���m�m*������H]�?�*�5m���z�ݾ�L��ۊ��ᘗ[��Q-��(�6�,FuH6���՟is?��߶�,k��[�G����IOG����
i�o��h��S��6j���␢?-�y�;*oλS���t���c�h�?������\��d�km94�I�Ļ�~p�>���n�sR�X��Ԗ2�ƽ�F���
0l�\=���K���R�ҭ�nE�O�D�R�kQ�/�~{�����-���|�I��_xK�k�δ3��$&e id�����&!���3�T����:��e�݄�T��2�}ޕ-�6���s�WP'T�m���)��c[�$8Vb�j��Ky�������\��2�C-*q���2k��Ͱw��,c`;�=��ۏ��M���t��C�$I��-zn� ����#J�.4Z��)�d����.��v�h�<�f��i^yK\I�P�Y����>fd��Q,�ht�.����jc�pd�u*�o3;+�~(|�ն�E����6�o�b�W�F��uh��ܸ+��hK����b�u�����y2V���Z������V���vMBV43;�; ��D*�7댯t�2�J�>�ţ�t�u3+��䒔�D����M:Y�`�z�Y�0<۪��O���Jg�ִ���1q��}W����V斌{�͛�JO�m��i���eZ
!{���/�l���VPW����W�< ���K���qW{�c��Hdf�zɠ(N�/�k�,�����YV��b���:��c9���o�{�Y��2�7(NO�<�6�vAy�e?�ﻋ2��.<Zz�x�y�P��;F�ɁN���wo�:�B%m���7�o��ݼ'���\�Qz��O���vw�2o{9��� ^7�^e��݂��Z;j)�M�vF�پ\IPt����F�u;���Yy{�\�ɧ0A�.;�i�d,�\S��%Plz��~��]>e���q��O�9�of��D��Ӝ��(ۙ�8��m2q�q.b@���cMyD0��?
��L�0�����:=� t_�c��� ���$u*����Ω�q"͓�W�^�g��������&yT#��}�{��k�y��SH#��S��UޯyK!��xΩ��`kww5&�N?�� t̻��i�}��졗����$�Xb9����*@a%�U6�!��;���;0�K��Nw �^��} �ne�ޫ��q@G�� ܵRm!X��]�
<��"!F���Q�zO���bfVCc ��>C`����� {�J���{�M�皐�U��v�U����Ct0 �	��{jq66z z�����a�6\W��ﱺ�5u�O���;�(d.�p�������0�,X��h}�9X�`�܇j:ZOML^&�N�	���������� ��:M���.��h��A�$���4�0{E�g^�j"hD� �(�KW��Zy	�Q�b����n�C�5y�2 �D�O�Kr"�@��^D�2彌@��:!��kk����7�^L`T���xP3����$��f�~��j�����1��ĕzM�-T0�TL��zC]�V��"V��g�u����`�=*E�!M�A��{��<�ę�!�"(IM��a�н���E��O��HqoJ)����v�|��te�i�aXo�2T�:�be3g=D�۴Jv�ۋ��P��_����k���'����j�����[�_a�Kߢ'n�'ߦ+%}�t���7ⳭھWz�߫3�8'�����c����X@�q7:�������4���sN
�~i��N��
�x{3�6>fΤ_.p6��)��#�,��V�op�.�y�4'��^�j2E'P�;[f���X��(5��V.}��pAN�|,�3uݖ ��0����V�6^��N����C��Ѳm_��e |"$�;_�Ϝr�'���d�w��.���.3T4c~���&��e����W�D��0S�I{��I�[��Re�'�*���!h�2�?����T�-sE��>L)A{֊���L��HY��դ�
�_�R�%dP,x�h�+�(���s|8O؉ӯ��Q��	I�L���H�כ�c�j-a�0����i�(_����Zz���H6����ּ��S>����3�����?�bOu�����"G���%��2X���o=�I!_-@BXOchX��yy�0ă2�Հ� Z�6��� �߫?b�.�nlfD�J���/?��G�+���2L|���-��Ԥ#�����ك���q�,��"Bj���\���Pc��I�ڻ�=����!z�y	�X,�LBQ��XBAR�|J|-`u��]"�(�e*w��m�0R�u���gJ>��q|���>h#|B�6}(H~Q�g3�a��#P�·�W�;�'�ȥ��Јϱ�/1�����ji-x�'�m�-]��mP5ҷ�T���H7����?�͘).�����#��I���hNTw�kMKwSX���s�5�gs�#�9�#��b��l�l�=7������}Qx�j�X�V�V��6E�}%�*�V�k�=E�m_d�v�XW�z��K�V�7����yŐn���ϓ����E�g����܂��&v��:-h���.������d�������RNZ&�nQgƪU�}��d�wm4�zs�[�L��ѝ׮�?#�/$���ל���m�{N�o��.���s ���yw���߀̺s�v8V���jy�!�g�+�(O�d���JC���x�u��R�����x�g��5�G����?+1|�z�A�D��u� ���b�O0�_�U��ì�a�7�3�E|��F��S�{�����
�饻��#?� ���Y�4�"+)Y+=0Nf��/�	�@��n�\��w� �n4�- �Z�D��}���U��)<_�]��KE�)���U�x�S�0V�c���!Qǵ6�V�1�rK��D��@���)ߴٽ�sG KF Q�ڼ7ZkE;�2��a,�"	*Ɨ����3�Z����c�=��bp���)�غ<��SX|͡��C,#L1��?щ�] 6�Y���6[��=������!.��E�� ��'�y�W��0k!�Z.��vu������	I$(V{����6l<��.�������S��ۉgr1"��R���&�� ��5|Ie1ɆU+�`����
����}�f�!J�9�OU�éhN�*1o@R'�eq�@����|>A9M*�m�t��+Z9D���0.���f�&TIaNt�m�EB[��Hå�C,�Ϩ�!��Oe��F�1���`�p>ޙJ�*���`�M��BP�z/�BE*��C�2��gdh���`9����|���M��U���1�+2g'�w.~�e:�xs��|��Oӧ.n��_����K�����:�6�g�*���(��<���^�~�=��-OitA�#�ZY��<\@>�gSڨ���b&*�*ϊ*ʘ��լ�-�`<�J�^������l?��Y���,���*�sfz:�����È��":A*g�׏Њ�q��wޫ�W���"�d�����/�51a!/~Q~er�S��;[�9���t)�1�Hq�{�,R�	���3��_ޯJ�yii��B�����\���-��vZxR�)t�R���t���ګ�dt�����xڻ�S�D��u�|ŝE�ty��rCϽb�?��N,���V([,�}̙�F�5���	��2��@l<�Lb	��<`�+(���4�z���'d��:V�Y�����^�aa���0���. �903��D� A����,�R�ۈ���6҇m"z�;.# �=e�?]��<�R@s�G�M�t��٥U��Jb��ԗc���0>-�RY10���ii��������2$��Xg���_^o�*�����B��F���y	�u;�V�	݌��<fբ�	�_zn���%)��{}:��J8'��Hu�3m(�b"�~�A�Y>8fU?��χ|��٬cR!��g"�$��� X 봡����0U����s�
���K���Z{��C�/O�j����Ni�<�R��Q�rM:ri�H\22��I�ew���� ����^����4�@ �`t��p�K�`W
����G_�H�&�^������������ޜ�RF�f9�'����G���]��}Xtgۮ�h����Q,x�2�+����F)�����t�W�"�;C�i�Y�����{��Q�哶Y3Mj>�0o��j�I�!HIi�͙��b�{fsZ�{������{���_�w>��utX�[VкkC6*Z��q F�=gf��+5;&\\�3������x�N|��W�bK]�ا���"��?��m rOy�=n��^R^|���������&�M���O�o550$T-dY+m�+�Ƹx�|����%#+��l ���Kg��!S��VFt�qU,0��]��<�A�ޞw�o�Nv��t.�.F-�4c��14������|���a:��pj�����m��4�!}��q#���F���+��u�uq&�#���������t��)}�٫v"�q]�` �:N�H��5�̚���	�bLP/�MRFЬ*�!CYQ��p����_�չ�y�@_��컻�8D/A�C�&�i���c{^�����P'�w���ú���a/a�nH���]�K ��u��ĭ��|j��2T¼�:Ʌa��l�5W�iIw;>�[��U��BFי���P�ZH�h��j�M%�[
lQhJ���|��B���,>���{:�w*��|Xa�x�:�����H����ɀ�}ׇ�:,h C9~<��B*},�o��{W�>�������.�����k�R�q�ݚ�q���'C��m
��b�6��CBh���]@�8m���Ba�Z������^#�R���^w��O%:tq6!]��4xg)1���H d�v�B���_�o�#h&؀w'sܥs�\CrrD��X���G�H��G�JG��Mֶ� zi��Ӂ���7�}�nhc�^�����S� �&X�N������F t�'��y�o��u$��j��~�����>y*u]n��G]t�X7.��c��ԳG��,H�:�� ���M������9�*�G�'����#2��W�|�ɏ;�_�8�^=o{y�y���{����%9[y��}9v͗=�7��5-�`eߏ)j芽s'[�Z��'���[�n��O�恾):l��|�Z�4�7U���a�cm��M�d�o-B�����ji���t{�F��/L�84ק���A,���ũj�~���gf�=�{U����_y�E>级�_��0frjћ�Oj�F/]��+k;7�JHp9}����kܣ3��,�'0��Sg�_�7[N'������8ȝq��/�'
����i�=lyI͈ �|�1vZ Q�*��w�k�z<���BT�;�>}U��c�*��0�x*�זf����uH��	̨��/����ǚQ���Hh>�oe�o1&`B~��QO��.���u0�pJ�9����Wc�Q�ߵ�r\'^��}E-M[Uit��]���[�_9��� '�������3A]�
G��-?TW���(ǁ*L�3"�1�f��20���t`� 	�ζq��Ax�Ε��:���=@�5~`�<�(��o��G��`��P�U��_z���ϗ8V|�=���:�"�Qv����?�$LbE�E��?�s{g،>���Lؿ��p�5��/�ϸ&��TYH��@�b-DJ�M��LG!G) 6�A�
� �����c��v3���k�L����\�Bih_<��	���Ɛݣ��YZ�]��>����%)픦Y� �8�.#sV��[���Y�in�z�ȱ��'9*��dZS�ڼ*�'/�HM�]]}H�����$<D~W� 29�k�>�/}�F�nl�%�H�,Y��=�|�}ݬƷ`��;�7߬m�|�?q�D�ޜD����j�O�=0���1O&
�	�)aeJ��0��D[H.�1�f�����G���b��u����^}d}����������Ak:��f	,���AM���_s��~P���a��d��gl8��� �ۅ�� X����g��Ԧ���^g)�s%2s{�ZH���l�e�2�e�D��d�<kؾ�]�ɺ"��4``��Z�0P��Q�~�H�X<Fo59���xD�����i`�&�e�˹&�� ��N着��E"�l��Y�.R��8J����*[zxF��[O��P��@�2gyPo����"���U����z��,�kͺ���$�)Ak�mB���q�Q�B��ڑ�6�6��R%"?B�Qs}8`�m."tT/��v����:+Z*���J�Y5ᣀXS� �������D���2�wE��xh�1_KRx���؟�b�C��5eܘ�5J²m s��X�4yˌ�i��=@¿>��:@	W|�����ZJ�v��zyߢ&��kY�r�4R�(�� �U�eP��32|���(���l�ܘ��X�0�lU*F�*S"�@e�1n�J�
���PF�7�9� ���7�1����)A4 P"�0����K�r¥we$i,c.�R�k?�k�8mQW:��tyaLI�JX6e�=FW ����e\��g�	w�Q�����`2Ȁ`��Lr�~r^R����(W���T���Lt��6�.I�"�, P
�Я+'�v ��c?��sr�5�kD��Nj!^�	B�	wn8���箂TF� @��������\�P�H[	��2̮=���k�J�X��V;���v���&ك��菂�#�Җe˷6T���d�YҼ���k?�	�u�ERK�d�<�'�q����?۞.�.��Y/� ���J���8�6�������H+�RV����ٮ�v�my�>6������cV6�6�����*��.�[7�n��g�J�ϲ�7۾���n�w~m��N#l]�vh̃��DjQ��P�ZP��;��+�:�?�:B@B�0^xxO���"CCl�*�}�Bbr�ĺ����Y��>{������ץ��m��ښG��d�KȪ��]���62$m��v-�,��@a�%�'�6����>�/{��*h��o�#Î��Ч��� �00u�F���t��<W;���g�`Dq��ڢ  ������>ҠS��s����6��B\;��q�Lx����>�V�S�P潻uN�Cρ}\��<)L�C�/6�J� ��C��PJ�r���1#Ɲ.�-�@($��1���ʹM�A90��EA�ϗ9F@��LZfyw�Q��ӗut�	�z��jH?@T��D������L�\o��Ae�q���"��Ī��G
�� ��t�цyKL�e�-	[	�༗�]��L p��<P=���q���.�v�*�T���!=����)�C A-U�<��q�d"��>��\ �W ��j 4L�!m� �m�RF�%��c4���W&�:��(������gD]w��;�>�r�k���8P���u��Pu�t-�7[�*�F �=}r����_�� ��X�>�I=�t,o�ێ�CJ��A
�P����L E����;���Vw\l($ƏP9���v�xľ{�3�_ޚh���^_�̾�w�`$��5鼵qv�M2ʤ*+�};�arl�L�Q�ź&]}�w�t�������o�����oh�T�����t�U���ҢV�Z}���J �#e��+�f�lu�A���3�N[^������i[F�e����b�bs��v��َ���>�>�����Z�l�~k��ϒ-YQ���/�d����39S��4Kꈱ��GV���˫A	 y���9H�E�u�
: 	0ᦋ@�SJH�:M�	j`��)�[��yH�!�B���kRH�e\v���c�{�;ߓ�]��z����{'�o�b�A���'�R�3�:Ǝ��cL	��qsC�:r`���0�h��C��$2�}	2/}��#�(a�ݭ&D'd<��R@�z�ἀ�z�/_���h �ב�|އ�(\+�IC]'��u&P�ך��Q]���ѳ@�q���x&4Pv7��k漴���"z���G]�?#�����8��P�@���y�
cJ@��%AH�����(��(1���xSݟAg�} e s� �q��v� 	�:�&������8�!H�6���u��:��p��H��p�1��H}2�����*����M�]Ʈ"|;r� �D0�/Ɣ"$�}��P9��W�11�$B 	��1)�}2�ԥO@F{�@*����,]�$` P�1#��XR@H ��(��Ε��`�Q'6�&s7�� ;�$��S��2'����!��t>��c=��ǵp�� 0���} '#鼬�$w�_�!�����J�./�;F�B��K$�� �I(e;`�r�8eƐ8�x�:WJRD$R%��� ׿WG���Yn�w�-�u�mu��|�-�?�6���:�) �k���U;�"�QFy�2�͔��yH�r��{y}]W����ۺ���M7=h'���-m�r�@��`)�������z�J)a��V��Vh���%�}�8�>�V�<���7�^�a�F��7Aw��{�����d����|f�{K��ϭ�@��i��F�RIdr��g9]�q���\]O�`9�������R5��<�K�Ϫ��f�l��U:���C�	�N����j��D� 250����r���T�6��=wٴ�_�(��RHSl�cRH�F�վR:���H����K������a8D�1��R"��}���#�r�x2�`��Fa`��k(�`�1�X(S�}n�(���Ĉ'�|�F�R�� �M}�80�@�6�Q�j�q^���JI�E;�UB�TK$��ýц>�Ͼ�V�s��B�������C��k&�(U����F� WJ�M}�֯����JP�c�>;�k2ڗu}��F_<d42?}%PyF�σ@J��Gd�C�g�8���?&>�~��c\�dV�l�� ��a_)�zp�)ʸ�8~E"CB�@	 �����_�vW���;���ޮL�V���#@� �Ft���>�Ҩ�;)�R�;J��H�wA#zoH�ʤ���nw��o���f� P�}�a��c��Xf�3��sF�>�'���,�R��G��N��(�e�F���Q� &/N�`_s��z{����FM�ȹJ�Zv侶l�'��=���%F]<h��;���R�e���Pn3�H����*�On�R'�����E�d�γ?�@p$6��M���*(�yQW�V�k��PJ �<ځ%�ܮ� g��>�����g����0����'���!P2cC��0�R=J�
�c���N@�8$cG�(٨���^�^���-�������->/�������-�zv{���� 	��?"�m��%�'�B*�E�<��&pZ(-α'��������n��ך�`a��?�v�Q�a��ڨ(3�=fF��di�+��#���u���/zo{*��ӯh�>�����X�^�����>����~��8�}q�/��o?0�T����`�y��v}@}S������;���y���0�5
(@*����	�4� qۙ�����d��>CC���R��Uc'����C:��k�@���C�즴�D!�X@�f��e�ⓟl��%�8�m�׳.h[O�!�U0�2��>��L���7�1fE��������Xל�xF�rػ�v�"C�h�T)	�b�'�Bu���&T����{پTl�J)�Z�
di�u(�Aכ�j�C��JlP�XX����C��l�i�^ F�~< �&�2�1�Kթ���q>u�x>�C�7��?��,��˽m�?��,m.[�q $1$���U%2���S�CŦ&��R�U��晹^�+fD!�B�R"�-/��k�9Ƙ�)mI?���f�=P�!��f *���-�N߬�כ�����Hl������k
�ԡ�d��s���r��z�]��O���$����Kt{������X�F�Dʠ�b�JOǠ>�k᮳ok�UyS�y[�}S�f(�$��1����M)(���{Jx�~RO�2?i����\s9f��3ƾ�C�+}���w�I6PG]�\ �p��(QN�<�f\�u]i�]A2�7�DUY)���pܧ�����2�e(
B�/
\���.�%�#�;�Yg� 
h�'W�:�u��@4&XYv�$���>�^��ۃg~�-?��vϱQL罻����kk΋j:lN{$����#���9�m<jz)�u�L��P������n\~:��vG��s��������9����x��q��{�!3�Oi�'���5P������m�<��:<��\�8�=mݜ��f�{�]������w�'�������7Mn�����ȥn\�vW��gs�{�s����w��$o?~^[v�m�{���;�����v��D9q��,�r�M($�h�'� �B�p�QE*�*2=�DIM��U��`��#1����}��	�ݔ���~�R�Ү�Э7�UbHQH�̻���������g��2��o�.����[�o %������x�c����B���|u��R���9O��+�I��GA|�;��h��a���C� �]��2h~A`J��j���r_�j@f(#�A\ǵuEF�s����+���<��.����q�q=)�R5�P5'�ku/�cG�ZI�С�jF�\�$��wY�P5�]�P_�RJ�R�978V�{����VC޼~�T�o����p��̵r�q�� �u��u���WًLX~?�,�g���.�$28t>��A�E�d܂�/QJ���M�${�&���k�/s���
�O�\���S�.=u��^gb�R��Ou(*��m˵Hl��Ȭc����+��k��ȵ����qJ�}�cJ�����*(�p�܌>0(����W)0%�=�t�SF���o���:���6*��囸JJm�"�d3��2�\ߘ�A(=���` �8��cp�HP �8V��������
iS�w�w��)��e{hR����xv̱g���������ں�������� 4��9zZ[ؔ�L�:H\wkA��:zv[�:+)�̾����C���}���oϼ��*Q���gF�@GG�;��=Jv݉mU�dn�55���y�33ܝs�?��rí=����9m�q���_��cm����E�0�m8��v��
8Wf߲c���.o7�rf�-��ꃦ�lKs��ϸ�]E)���nY y��BS*����P:�T�	VŐ*�!�.� e�eő�R�yҾŐ~~�����ܓ�|��5�;xo��;_i?���~�����l�,�����?k��wY{m�e�_O���6����ܷV�W14�e�y��{��%30H2� ��R�3� 0��8����Tj#��>F���"�)0�i㮎} d�N�S$�PKp�8��8n����R���,�6��|��}̑{ �:��� �k�r�����7ڈ9�<ʕ��);�_��|r����3�� "`"	�@��#�}7正z@Iq����B	ؔ��Җ���K�'9�Py�U�|��!�"�A����[�c0�q5j`��Z����r���8`Q�sWC���V�vi;�%����u��k���4C*a�(#*�r�bH5KD����V��:�('7���PN���<e1���e�N�T��*�#ޡ�>sԊL���v��9�8V�so�6���`Z�Î<[)��w5���p�(�2�)�H����n����߀R�)�$�q��(Qi�Qx����9u_��! �£��4*��+u�� 6{�@�@,�U�Rڥ�:�B� N�!�1F�B�e+^�z��U�C�<�~6ƈ���@a}��-�g��G�^����W�G?���Yom7ͽ�=�ϵ��~�V�8�-Ir~+��:6:rZ�#n;j�|vkc����Som�\���[����?~�m
��|�/��������= ��1_���m͑� �Vd��������m)��40]>��v׌����7r����)�_����<�y��%��%���/m��[g�ۮ�8����Y�l��{W[:��v[~�u�/iK�]��(�b?o�u�z��8�\�,�%�e���� ��AbHc>;�!���R 	�ј��d��|�I���.;i�_�_i_:��RH����+���H{�n��-�TR���Y��W� ��:����w�eS埕1�� ��=��3��Ҭ*�zg�y��uΥ��2�tŇ2��ؗ�Q��G�po)3|�I�`,{�i��RRV�1�>o]w��	��SFދ'r����票����B(���	��p�J��N�c�àHlosF�]�듐�ߝW ������'��	J��HR���0�)STmr]��ӿ)�%e�+`��o���ݷ����y����>s~O�E�p]My!H�S.`�Rc.�!�#P)��`���q RGbeE	U9}t(M��R$>(Sd\~[�F�7 Il0���.n:���]u���z�d�C��-ǥ7�@QWc><���S�_��6\x��0�"��<`3* �X�x~0�#ܱ��O?�T�R��E��<�  ����K��Z�XT2D�X�d��RS��(7[��k(��R'��c�����s�r��@4T��@���a�ws�QJ�2�@��N/����'QI 4�P��#{
8��Cib��R�/=��Cz /R���j*�=������^��O�+_�N�o��E���\��Թ/�K���4=p�V
I2���7����9��͵�I}3'��3_8�vSѢ��U�_X��Z�c�>5`1�*etR�7��>"j䐓��(�I!�s��� )��{&罻=q���#�}��퇞�<�����h�9���Ok�s��ͻ�����mi@u՛����|O�vŧڊ9���~wŕ�̾�/�h[�N7�~�L��,�W PꮺEU��:����($@��J�TŔ�J���7�)]sP�dLR� ]yȤ	 ��v�)��p�ew����7����v��׷e��t{��K۫gG%�>��<嬶g~T���1�]���#�h�LIt �e�9�,�aL#����S6�:��]|JʿN��`�?��M�)p`P�*����}����ư�0 ú#�L��ñ��$` ������s�a���CΣ�kWǵ�O�Ch_2����Q��6�?�"�N�p���.oH 2�s�5���� F\��d�pu�wK_2뤄kT��8�g�����d�X����$yEz���ku���ve`Ptx�9H��TP�]�7%%��l\r�bB�;.����̥�x�-τ�N��B�3 Ҙ��bJ�n �vV}�9'.D)نNL�*�;J�PO�H�S}�- ��o��s-R�M�
*&;s��b�\�()�%~@�����ۡ$�� ˕��>%5E��RI��L��_P��@��>�	,�J]��1 �FP�I��g����\�:~`����X6p*p�R �]��oʠ�>�(%�O��pՁK�)e0�*�>9��,KQ �Hh�i���G�
d��cC�N������Ҷ~�����E�p�US/m��7��ȹ����돊�82���|Jk-9A-1�y�+�F�D-�얦��{b7n�3[���y�K�Eu�ٽ�I�������ޣ���2��6�:V����e�cq�aӻ>�v|��ۓ},*�����s�/�[z��m͹o+ �m��/i��zv�+
��(��G�mw�nȳ�;��=��o>�ݒ�&�n�oqK`~��S��cg���4�� 4��e���D����� FHbH �/��W���o<��nc���C�r �7'��~�1�}���'���^س�=x�Mmŧ?�:�.o���Ҷcz�9��m{���b�To����$:�R�Y5�W��8丷�W�E�DI9ft?�D-1n���c�)�� �EE�~�?$����q%F��d�A�qT���a����>��7�,�97�S�rL<�����N������(9j�_k�e���V\�6e��P��ݻ�y��z+�#��r/ ÕJ�56#�T1��OL���1�Wc��,�ft8�+�\c������\��I�P;���۔��o�(�o�A��P�(*G\GJ�$�>]i���K`@J�d6ѓ��J9��B�T)��>ԧ�d߁`-��~S�JbH��P8J��<vy9ȳ5v��z��������PJR�1ʳ��);�N 2P����V�1�
��sw�~A㱜pԑ�`�Q��}o)QS��r/�g���}�%#i��Q~pĈ��l�'vN��R����f�@K�+I!��m  m� F�rץ@�*����d��Z�bN	�j�캊!Ű�����&T�p��b8�ƌ���_�Ǩ�r��>��}9>f��/ꣀ��6]��������5����mm��絻g^�^��ּp�<"�����!}�L;@*(��[5v���\��\�� `I@�"�L�[�����{?�����8�+rNYr}-$n�����hĕ�2�6R���(Z���G�Y�KO��ݘ���C洕'������چ��n(��WG	������ծK?�_ؖ��3����,��zdƥ��<˛�w�<���Fw��-�2�9��=���W�3�
Hwp�������9��xѱ��j��C;�*�D9EI]u���'Պ��yR�����(��_�4���i���[�+� ���=v�¶�S�����Y���ο��<�¶uf���3��b�)1���Hb��,�8>�(YʼfH=���Z6�_�o``���YƑ�6�v��r��K����ql���`�ry�p1������q�,1�h6���b�b�J�O��_� �:m�)�=F�r��\;p��6�<�k��w^}���j0Lר,�Nv�i� �;�rRV�W���H
b�Nק\�$�Բ���q]�\�X�O��L(�W�[��w�g�s�h6��ʒ�A.�(e�;']�]O�>?//�}ռm���P��J�q$�"J����b�K)���UMW@fh���e�+��P9 "��*�T��������H���(���0�bG�hd`Žg���7Ԕ�f7	��]vSɔ��2��՗�H���)%㭍:#���?��S�+֓��� %��r+�J��@dۙH�4�� �O��#�_ז>)1�я��:��،?����8�;(+���򬴫	U)�|�Lc)sЪi��[��T�(��"u�*c��g=�Gs�Gr�����ƃi�1���t�/G�����������vÜ����՟��/�H{����1��|j{:�����#I5�ݡSښC��5���)�<jV�+��T�|�/��s���;���(�3�=y&G]r��CZ̴��U��̽�� �P@ilL�X������o�d�=�+783�|�zO{ �Z6��vC�W�翧�{�ڊ3.k7f��g����z~{d�;ۓoy�-�ɖK�O���Ŧ����ۢ�ܜ��n?lZ[ K\��H.<�'Dq�;�`�eד�owDMʬ�1�y�n�l9�]��9����v��jWrl��/��7�/~b�����|�#��������v���=vע(�?m���ζ'�赹yc�}n{e�%��S��?L�1zt�Ao�S����l�wU���[Ŝb��qo�R�vFJ��Q-�2%�N��0� "�+�;��p�Q5��21��g�s�u��cJe�sM��P�bHٯ����f����ڀ�rP3��0ڮ�!w�U'�0�@,��1.1}��>�\�d����<ѦZ��kC�(0�ϱ�p~; �ֵ;Ǩ��Q�c�:/~o1$P�<�l{g�,E<�S)�y��F���.
��m�
X~}�a�V�z��Pc���ٛ�7��|)Ywf�3~��-1�`2�L@!�| ŧ��M���/
i(#�Q�/�Pg�un���l�5�Z@�1禣�(e�^R��_��ᮣ� H{�!�����`��b?��S�{��2wY���1�C�>H�/xp�����N�9�G?�9�6 �O𡂜�
s���<ʀc���A99W�o��C�9)&���|>�~�S@��&�Jm��+�R��� �m7�=���e����9����?o�����gs/mO��?����v�[.k�����;�}m%�_@(<���1H����(������Ī������ҏ��>�'m�e�o����m�>���^��
Z�,?���Ѻ��N\u'�:��ԁ$��}`��Y���G.�X{芏��s.)��ó�h�H_��ȥ1�y&�b~��G���8Bh��;��}�a����y���xF{�⏴G/�h�6P�&�)�7_��O��S�j7�s����p;��E��>j���Z��2�!ʈ"���$P⾫A��J7��5����_D)җ�8��ŉS��?��v����~�e�s�����w��������n/̏ژ���=���y�N��+:��5戁�����F)�qH�ܡD�E�Đġ$:�U�(b4���5���PZ?�w��� F�KLX�]�:T	��>�N��7��z�<�����1���PA� ����>}2���W�Rw�����
E���;�����T���=#Yp�z̵�p�T^���q���\���{���Kܪ\m������\���>dn�?����L� qY:����(�K*�P0@3�A)�W�}��b�z��"^I1� ��Z�/,��UJ���Q�ڀR� )��v�p�v�<C K�s�Q9>_���ۈ)s�HHI~;���#M-�d��
�s�֕R�*XJ��Ў�$'PA����"q$�J��wj��] �r�K?���*�V�� x���3p K��p��?\��\��ҿ��.@��1 �~�/�_�
t �~ҿs;^�&@5@h�Vue��֚�!�k%ڂ�)@�w�?�}d�R��5�(P��:4�9(���FI�N-�ύү������Ӷ���^��Oێ/�=��?o����m�]��v��3�=GNo��*���c�a⪛�Ϩ�cf�����cm�j���w�=��������������w}���o�,�wo��ܲCN���J����|r[vP���F�h�����|.�v<�m�'���?�v[���o����8��s��mel�QX��wZv����-]pY���QByix���|�-�rV�q h�G��G����8]��_��f��ɋ>�V �!�=2C�P�LRϮ#�:�͇��,CA	�Hb�)�h]et}��1O�T���?, ���������B�E!-������
H/�uY{���a�m��y��s�����K����,CA��y���0 D�X�@=��i1`�B\w޶��u�\1����V��zJ�Pepc\�QfXGV������0�`@U�L9TI
��Y0���[	�=��!�p��S���� ӨC�T9}��,�y��Fpp.JI=1+ t/��������m�J���.��}��5Y�1�:�ˠ[���y��Z���:T����г������y��9�}���3P9bH@R��|�ŀ�Pɾ㾣��&m��� �L����R�-u).�;.?籔����A2����kR�{$6�̹1樻��nO�Q��~u����3ؕ�} ����ԓ!d�Y��)G�PB��؃K�!�x%���]O��㔴��Zٕ�B��Z�9�x3���C�2�ԆX�ą�X�,
J��e��z&@UG��F�I��2 b���9���α�N�T�F�RA�G�d�#u�$T8���f	�~��Kp $p%�Q�բ~}h'>�D^j~���E�d�9�!�ۘ�7�9?s��ێ��v������>�����|�m��o��?��mټ��]ǞVi�b7뎘Ziޏ?��[ce��Z֪��6׸������>��Q#�n�x�᧵�d����Ʈ���� ��aPEaq�D��PL�� �v����Co}G[2�����jw�ؽ��8��m�������r�^���]�w����������k�.x[{�����������Smɜ��C�}��;�m������6��wy�9 ���i�<��GN	 �o���.�d� *�?8�]��c�5g��*�TJ5&)�\uD!]c`�Ƕ��A��QS�_�tJ���>�n����U?��B
�V|�s���^���ٗ��ϼ�m��ĩg���j��3~���Rnh*�;��95�%��ڗX��j�Ѧ�U��z޾�
�b@cD�Oo���p��pȧ���H��PB�kWPʵ�İ�$T��5Ȋ�F=�J�������Re�<�PP*������� ����>r�����< ����E�cS��ܓ�q��&J)���k�rY����{();��TC���k��ԡ�(!���SM4����-P�����]�]����r�A���{Z��c���S/�p��~�$���R���Ͻ� L���LI����"Г��31jCʹ)��bLM�Z�y��pí(R�G���	`���ϳ�1��
0������S�������$BPH �\��le���d�jPR.�X�BJڨC)�-�e�2�u���PB 0L)��/����=��6 V��	HY�t��k) z��N�Qv�zK]Ɵ���9����� F��࣮2�q��S�J�`¥�f5�CT���Tq�x:�f�JC*����ۣ�ϋЃ)�D��1�ȵm��<p�m��w�U3���qi�#���[n����4�u]�s㡧���,��1�2�j��(�{��mC�I�0iE�}Y���Ɍ�䚗D�u|VI�H�e$\�H�����7TRWG�}I+�ЖN�3��������;����)muߚ��ێ=��=�v{ο>�]�����w���/n�K9?�����0?ЖEQ����me�Ć���=t�{ے��\�g��̀�ҏ�{�~W�5���)�C���"
XF��r��L;n: �)�T�u��{AhJ e��� �bb�/��
H~Ҍ���},
��QH���v��ڞ\rw[��?kO��}�3��Q�F����[�~=�S�u��p�>��)ێbb� �*�Ę��j�eʔ�2(1����SJ�@򏽿��1�յ�q���>�M�~�
��cX�X�1f��
��ap�����<̀�ր����hc��H�ԉ��m������꾄F�i{������Ղa�	{��9�����Ɠ�'��y��9ܭ~[�$h��~�+���^��;.H�,%�0P)�@i ������=�>A	�F�}7��J�N�gcȴw������{���<_��ns��m (�)�9		=�����=��]o�0� ��cF=����r����q&˝s�=�c?���?�D���Sί�i�� �O�e��rO 5fx�F� 3� P*'��>P2�R��E�Sb��)P�ljPk�[���-W�sҀR%P��
^q)�N�*}ed�M-��7�s�y���|JtЎ*Rvm�T�¡Q'y���cH3*�a�$@*55%�z����-=x���P��)�s�������ϴ�����̥�n;���E�h���_h�μ��p�vH���i��eε���IZ-�e��Z�M֞�kr�`ڵ�[+�xV1�-�B[�����fVj�6LJ汫��6pꮺ��:�l����@i�9��g��S�U��j����2Zuʂvϔ��ʨ��s�˦.(HY�|Q�rc �r�9��h��tF[8iN�1�t�Q��;b��|f�:ױ.jk���lO��my��V�]�W�m�ʢ|.�&�� ���W�7����w��8�Ϋ�p.�@궨(@���s�c�Ծ��Ծt���'�h?����MQH?�Y��}�����%mŧ>מ|��ۋ.m{f�`��?�Q5s/j���Q��=(��9�c��o('n=�;u*�#Wj*}h#�$���SJ���x`P�b�h������r�n<��㎔v�)�L@ȧ:���P,;�s�ʙ��>zF�F٧>�)�aλW]��}3It��� =�Գ���6���.Yp�Z���~��kI�W�w��p��ۖ\n:c���`i
�ݍkܔ</�ٲ����P�\=���
��M��p`޺���KG�p�� �!F!��G)QN�x�!�.m�S�)}hB��i�z�1����ƚK���K�<�w�X�\�P��W�vf`�m��QJI{)���H#�a�kF��P����|��=SNc �r��qJH�]�+up09f���]˅������@G<c�)�Pr�>���JPp��r�u@Q�K�P��hu��`���{е:רZ{�R���`�9@���ﱒ�fd��R���o�s��}c A=��G�/�Һ�������~�m����/}�����m��\[��9s�=��� �ɨ�fۘ��6PI��:F~��S���܂9���us�1Q�r�Zy����:�SH��k�m�ˮ�딧�옵�N�E��0��r��v��9ߌ�2�/5�'�;�0���6״4�f��[��8`�+����ﶜ��lw3�ݒz�M�Ѯ<tr[z�[�}翧�~v�a���GN)U�0����a�327t|�E�֣�����*u�ȮS����L�R��u�N��XK��������K����rj��'?�n��ەWRH;��gW,k+?��ӗ|����w�B�<5o�ӯ��&��3\;TM)�jo�� ð�O����mG)5�������a`����%@`�ap�lm���!��ZJ)�aH�q���b����2�6�E礞\�:�}�_Vp�����s����':pŕjK�r%�XJB��v�c��~��zpp^p�X�Ƣ}ڌ�r���J9/e�'���p���<#s�m���r����*�뚞�p~}:�k"��]
�u��aLԡ��"e�F�6�HbB����Լ@D�=�'\��J1��6Z�N�H)�U��5�Đ�ʵ�<v���R�,���|M�<�%�GY<�|�������QX��P`����;�=cň�	e4һ�R���bH��v�7��$��6�y��ǭ��&f4��s(��I�w@�̾���/xPL����oJ}�*�[�O҂>]Ø����w��ܜH������;Pr>������Uڀ���:wڍ���Ŕ��w��YRϽ �����_�:񣍇�0:L��5ݛ�{���m�_~��h��m�G���˷�i��x�-���<����>�k �Ղ�����Q;kr^�8<���/�^��r��nk<9Pw�=7�&`]e�:����X5�R����:nnAh���'\z3'�N\x}�ɒ���\֞��me�R�ʹ�hwF]�ŊCNn������m�RǦ�=i7�%��4�U<(P�9�kù�l�{w���9� � ��hQ �Ж�{W����/�Cq�]��G�Jc��+(����3N	�=>}�X��8@�����W'Mo��ݏ}�]��oM i�ֶiՊ�*@z��W�7gƸ�`�O9��k�K����6#^D��n�Q)���޴Ō*��?|���h�/<F;�5�P��	�M�0�ee��;c^��cp�m=�+3��Ne���z{3���(�_��ٴ� ������ J��r�����m@A}T�y>��׾��I�<u���ka���<ڎk�x\;����q#�����bq� ��P6����4CcƇ��:~�M��z�x�"�9׶�ze���d�u��E$e/�f�O�c�ە�-�Vb�" FR���gu�]��P9\{�����ȵ���y�
l�����/��!�u`�)�+�� �gԳ�r�闢鱞<����F��瓻�^��{϶�=�>R����R@CQ_��x*��qH��t�]Α� SƝ�NbC�����Ԑ��6@�1(��� �a�S.�W�`��( ���������q�pP
��>�t]�\��5�P�M������r�q̹�2�Y���\P� �~�|�?���:�>��3��S���iSO����}QJ��H�罹��>�Wm�������?n~�m���V_�Ѷ�w�e��V���x��m�U#~$�lҗ���G�Uc�����(nμ�Ⱥl#��Yzbu��6*�2�����m�m�!�P���Q��Ui����9��g]Ҟ��=mqε*�'mJ!�tj[#�t`TU@���9�ӺK�
L�ڲ\�=�ҜcIα8�u[ x�1����.m�O���z�i�[k�)�:��B���v�D)l=��؞�}�q��}QE���ٮ���������?��7��7�bH�����?�v��Ͽ ���6�]UYv�i�=����y{?��91tSb��OŨ1��$�&�dց�$�T1%@	,ď��:#�R�dS��8�?��$G0�e�ӎwN��AV�kLN�PW�(w�_�c�K}�g���t0Ӧ��~��5h�8C<࠿a��{�'�\��m@�f��_�߆��2E��V:�(�A$%�$C�rHw���#F�tMJ`�Ԩ�t�x�>?�?��s���~�|���ǎc�(��Oßˉ�uܖxߪK����*̉����O�sX�?�a��&G���!��9��(}�Ie�'�1�:98������#~��ձ�</K�-��O�A���a���κ�R��t�(%}%A�n;!�:j�:
y�5,�=ΔњGH��l	y4�"2�7
qxB����jq7Ze�ZfFsF�m��/m\� -����������+(;��z�lHk���~���n����n����TGge�U��?:	)A
1 ���v����!Ѫ�:v�G�l��'Ѵ�9R�T�0#	3./i��ٰf�7&|P;��rL���#�,q�)&�X��)�
���m�	�4�r62!����kF�HZ X���Nm dd���MF�����4��+ͧ��*�+N�k�������趣�j��m[Y�I�^��җ�su��G��r��鏊����4j�ꓯ,�؜�(��[��Ճ�`[����v��ZE�Ǳ������}��{��s��|:�u�}S/B��K,s"&������A�=}��히��X�&}�@��|T"L�r}�h�K����VǷx@�6��A��3c9h@S&?�"r��n.�ݖ9�a�d���>v��~x�εЂ������Y����u�� E�o9cJ���~�T�[�9��r��-8����&.�#��\��.N��d�OI�'�Z�S5^"��r����/����3C�
Y�D��<o\�BiW��:����~|��~{V�k'E}S؞��+�DSWgz��]M�~˫˘6z��c�S�Z%J�C(8:��5k7����fp��L��\�J��{���UN�bO��W�҇g>�և9W����n���kt��|��HKQ{\�P'�}&�m�����D�X0TFj�8a�(��((�خx~6-�UA��ռ�f�	ψ�3/E#��d���c���+����kc/4g�}N�f)��w��4 �)��/�#�w޻�җIj<ᒷ��Y#�$f��":��sm��b����z�oZx'
��}2Lݵ���������% lv���:(>���FU�z<lOh�����9�'���Se��W����+8��G�\���fv���(:��n�ʲ�C��T�XrT����;����a���0Z����
'�m�pZ*���4���~#��� ��a��̟̃�aA`��z�H�ʱ�P��}�#�3n�)��6���G��	*ij�}n�74�.+�#�����G6��l���0��v�OAS�N?����?�_��m&���G��Tfd����#Eܒ��\���4�W����>ή��/��#G)�r��S��Tz0�[�^z7ij�_� �� �,�U�-�;5@�;�|_�m+l�� �k��n���7}K�5.����������Q���m��r�r�@>^f�{n�Z��#HQ�����RTr78�B+���+�o.MeG�Uem�cY&1c��p��}�%�~eKrM���j_�=��H����o��RC���3dK�e�G�*H*E�D�^���I�~��=qy:X_�$��_�a.��:
��;�c2���^�k<�ba�x�m<��߾�l���H�T�R-+v?�-=��>	���=��oTby ��|��{1�ߋs��o�oDKr!ض���������}� ?֤[�|��%���J&G5��17Ǩ�=��F�_�My��&M���� c���Mgg����o���/uRJ#&����փ+��W�uۀzS����� �c����E��Äq�ذI�������f�s	V��!}z4��(.q��ϖL���6�k[i��N�����`K�,��W���C����LK��#l��_;7��-���Z�D��5��n�q*[�1z��	�{1J1Ю�P3�$j�GH&�8�_Z0��롒��j�u���W�?H�z��O�L�~\d��+�!vD0��[������u�,f�ǼN�`��~�
R�4���n����e�'��2n�g��yC���=��!��'��S���z�=Ef��q�i���3�TC��5~��T��.��W�.U�*�F��������yQrd��:ѓy�	� n�NI�d�6�;��9��N�� |"�*���wz���;1e���ޛ�#C�E��|X+�`�<��͛˓;{c�?�����q.�D�ôrδʙ4���TbK�j��M���-۸��n0e�������g��&|��}�S��� qST���B���ɥE�ly��q�D��K~��Vm~{1%{E���]�v7̬�s~����v�@$
+U�uu�w���#Ay��/�W�X��)�d��k�6m��1���w��c��msy���Ox�،'��*�n��Ku�izS�ko~�?�gR@Qa�}O���@V1��У��)N�J�[ϭ�7�N{������ab��:��q���)��a~˕x*�6�z�G,y.)�L��������a��E��a�Ʀ�׏��lכ�!nރ��+?E]~L�i���,[��C4�:��`&Hc}Ef��&齆D��Hg9�=%�_�<��T�C>F*�@��m-��WM��Ծ6�܅�I<h�8㌱�t���<�` �٫���x���L�������R�DtŜ.���KS'�RW��[��J��@Ł.O%�ԊҬ[��_�lU����@�]J�f$�d�ܿ��JJX��}~;B\����b�'#�˟,���\���*�>s�����W�W����,r7˄y�f���eH(��Dy"��?r����ù��	�S�o���Y3��4��L%����(�\)�P!6|���	�#��jf�Q�7!6
+?&>��Z
'oXV���:0
"'����B�p9&-`����,l�	wr���|�?�w�fl��0����팆������P�Cj��tzl(���0�&����lw�)H}��ƫ�*��ݠE�e�X�*X
���^����vFo������sks��F�,���x�9�����~�fͫ���t=�UG���YO#��3�;�4�������� �m����y�'��s�rf�{��=���V�z��fդ:e6��_�$���1Ebc�����πc{������K.H���ϸ;�:��>��m��[O��]�Bb�)J�6��G]��s����Θ����qCvy���ܽ�A�y�-���a�����%�տ���4�54����D���?�������k�	�\>��M��x��A��Z���G%��M4a�Q)%�����B��O:�3��P��q��Jm<�e�]G��s�'�1F�� �v�=��W����~)�yT���.�v!0��D=7��6Uw��~aT��9����:1������}���<{%��
6#{#6tVᝫ_�VQ�Qs���!��ǂ�l�	��[\uܨs��e2��o�
}`ad_�oX�j���~����qvF�D|yp�[>>󑁞��LF��׺�Y՟oW��v$�쎨9���	�
31c�Y��P�x�G?���ы��	��uw�f1�أ�Hl��re�豔�.9��'��,vYc�����	������{A�v�sm�Y�S�ϣ�v�#���������Z��T�if��Ev�����R `���-���D��|{��+�9P��o���U��9��O�)��=^@"V��k\�A�X��UAVKj|��L�ae���>解[�`�^{�
����B݆����|@��I�!�L��ӰO�a�(<2�����i�Ǭݼ�7�]��3�/ �
�tx� t �UqM@�C���ח����I�x�$�&W�M|�4~x	T��'I>�S+tPg�۫��;Ľ7y�=��`��qǡ����ǼhI���fU�`u���j:�ʰ�I��I/�w����?���-���{��IY�pQ�@�o��4/�m�w�c���o�B�\�{*'P��ab��������+|��wX�z�Xd�!
��<�2��.Yb�۫H}A�Ϭ�<ϭz��-E���a�멛��ݾ2�b��M�|�p�;��&��<��Faɓ�>����L�߁j��L~��ǉ�}ڛ�'��Zm����KN=ׁ�x��a�k������q+{��[x��:�zbT�M����{wrOk XK��+�!��$�L�)H`� ��������ڃFI<E��~CB��O.���!�P��v��ῥw����Ǎ��C�-�3S|��n��>�E��Ę{3��9�:� S!+Ҳ���{,�erI�JyY_���p�8�l�%Z�����q��7�ܣ�Ll�p�B���Ȃ��z~����Ni|7��3ѥe��g�,�f�i��w���0e:��[&>��97�#�z�`�IL��~�q��P4����&���v,p+�p���X�J�����R�{�a��r#�,�{�;;-�فR>Vu	��6�q|�z���>}�F�Up-"��QѰ/��r���:��<,�*���E�{�#�Bh�1�E�5Z*˽/�#�[�����6����[��E7v���wX�7�$~O<�4)SҬZ�<ϓZ�����.�v�)߮�t�W�%R�H$H���;v~ܹ���QSLs�1Fm��M{�줌�x�0p�{�-��7PrbP7:�y/UxT5��;Z�J��L�L�[�ϮWgْ<xM�E�@u�!�T����M�h��8�TG�Q괝t���?�G�e��R�T�VFE�����@H �R/&$�%'��O\gE
�t
� ��>��؍��n ������vR�]�fU��=��E�_��et�Ԑc�[>��H�cn9�*��]��CeH��ߔ��b��jqM?�lPu��37}t>9����3���,#)IQ|#n�\���r�^�^�������b�-�ǒ[�ЂzC�a��ס�\����ĠZ`R��N�\��(�/�`Ia��n�y3���%=�~<�.8��l���A�5$���x�`��D}?s1I	 �UĊ>R���g����~�����?�A�%�K·us�����]��ι�i��(�7�͘�Ő\�F��26t�O��@�'�;�"��/�'nq4r�x`��6�m�la��;n����3u/U�l�${�t���aɹA5W��b���s�KX�J�Bi�x_��6Uw]<����	\m�3��|�*�C�����o��G�=M�7#�ͬd�|�B=Wۅ޴6H��2�#�K�l/�%�� ��{�uuz��t���/&4�b!��`�^���*���P!��K#�R�}g=�Q�� 0Vu��R�c���{Jɟ��+
���T���
�@��i�qv�&XN%������0rbw6�B�xڑ�ߊT���.=�H�9�T���@$�#���Smce�����7�n��s���BjK?���D�?L_gᣍ�`@ޤ8O���R=��e��(h�_��?���VG��zly���}h����_���+�ac9PD���q�jw����X�1�a�6R��nѯ�Cc)�q��ޙ��B� n��J�O)�v�r�t�ǈm��Xx�4mB݆����]Y"qȫ�LE����J����ݏ-*͝.Vg� ��P�
^�o���a��(�R)^ �ꝠnK�6l�B��C6�H"w��{��4�.َpiڬ�$އx�qU��	8�:4?�����/�]X4�_s��}V���?�I��ֲ���r�C�e��Y0�s��ol��Ę����ʋtN�R!^zR�=+%��f0 ��� lv�b6��l�v3����@W#��Lo+[딪ZĔ�u��n?��v?��ײu��^U���EqXm������	�"�Y�Ž��
^j��m��O�E�3���Poy^�p]���m�St����9|O��vl)��������ZI�HQ��j��/c`���� ܓ	�3�*H� fT�$��x���'�@�^/#a:S��i�����[_8^"�cs��/������ƽ8jb������gu؆r��u���.>2N*�)h�ҕ�m.0M��\��@�u���_�'$���5r�vU������d�"�M��\�6ާ�,�� �l���M�+Nʎ	��w !�U�Z���j��E^��o(��I���z����o���&o����&o>��"�H��H�/x�ɰSb{��y�#�y���[���1���i�˃5(��?�e[�5�"��Aon�/���R��������m⏿��o�y>���=���ַ���K��G_��͡k�	5�γ�
��5N�LI�jX��]ە�ET]R5��t��Wg�>x򡜢�Y���9ԡ�����ѣ��GN���8��иoB�+� >GU��]Ap��Qp����,\�x dy��`���I�o0�����0�#ca¬�?W���Jml��O��0e��S&�t���E�խ���ҧ���S 7�a:�H5=�X��P�b�1�oڻk��`�-�Wt��.�%���/x)`*=�	���	[��Nc#Pr����8�N��w�U����y�N�6MM����s�>��)����lCQ^e���S��8b��4S�R)ض����O����F�h�,��_۱7�&��z�XZ"	K�K������޻��t\=wk�rŁ�*��2´��VI�� cӔ'T�1�7J��Y�GC�T��ݹ�]��;�͍$[��kx.?�w[��j�rC(���Or��y(����}��u���A���+W�'%벁_E�gӹlz��D���$����=���u��ZT��}�)����q��?��Ř���]���u#9��,�Y)��p�x뫧�����ڏzkNQ���Q���1�G��#�	���I�'�J����[�ǺGFl��E�d�a�缒�����e>R6�L�,/���b3{����ޡ�T���m�9�B�J�p��t��s�m
�4��.>y� �~r�����Ӆ��
.�ӕ��xn��%���_�I��0գC6G��,]������� މ[ӈ�	Sz�������T����H��QU�鑉�O}��i����V�C�qz:��5�C��~���)�P��ae:�����O���s���*��{�@����<��W3�����+� @��Ə��j��9Irg�
�}�.��2�
�{�"s�M�\20�m7Xk�dM���b��
�'��U�E��{)[�k�����) �v�XI��0B#DCK�R��4~��^�!t��m�����l �hMr'ø�1�	9��n`�νŉ�*=��ϡ����j4>y�9��
���]u��S
����!Т�A�Ϋ{�>�������>'2�e��B2��3�0{é���I3B��Y��
ک���^��(#1�Qz���$�(��Ҳ��.9U�q߇�M�&L�ӛ!���xh,���<1�"�����1��5���2�t]nG1Ҩ��Q���拢�A��D+2bk_���\�i0o�׷<�̈́ƈ�@�?��v�O�6�۟���"���/�=�"/�����ǹ!�"O&�溨���U�I��Y��|Q�s�Pke,���m	�1���W��'��ʰ�Ӧ�*����>ā��hzEs�{��M�5h���-�(:tQ��4�����;Ws��BEH|y��
>Ӌ���]�.�~c)u��m�z	o&�ZU)e��'���l7��z�����Ղ��~���YK�g�}��X�m���j��\�(�� ?51�t}�ed �<��i�
U�W1|Ķ��[�IjnJ%܏���9zy��=֮�A�qA�G��వ��nl�)Yv�ƫ|��9�7��91ų_����[�0�.������9����I��g�	�K��>�U�q�h�J΂�=q�����0�9Z�yBWq�@���������6�Mٞ���)p�]iP��]��v*J�Q����sa:��3 ]Ŭ�<����՜؛�Y*�;�xU��tS���󒭬4M=���wЌT��qy�kC'(FG[1���o�a
z���2R��4���Fܜ��6Y�?�$��ŏ1v��ޕD�BnN��&�|��z�� xLa�wx�h��'�"�]0����]b1AY��a����a��V���M�=<x�	jR�\e�tˇ��C&wG��#��pb��_��E���I�������B�p�yjs��<��������� G���(}�#DQ<�:A�5jXYO-�F�3�4�r2rM��{�M��O{�P����>�R���U��
 ��$if�޾�0���b�1�W��Hn��H�a�#R���ALC�rUE�ߗ�����݂���cP��\���u���U��9�S|���u�����gT��zI��W����Vs����HMrzǥ3�"��������~�pD(���"7zyt\�0��Xgm�ܹ4[�Pu��o�u��(�V��Q5��;X]���6��%��E�18|_��.x�*`<k�I*�U|�9V�`�?�ݸ�n<S�a�:��3������9�GA���DP&��M���y�i�U��
��N��D��.Fz~^&'T�y����X��	���ë-ܴ��驏8X ����ۃ�
�q�q1o��s����h���y6��#�i�̈�/��xW0�O���%5z8N��D�R�0���ǘ?�?��?O$�n	�@ʫǉ������v��ey�����%����l�(�<Q�O�}�(�Ԩx�Q���9�p����O�8%��Z[���ŭ�+\���t�4�l����D$c0�\ֲ^l���򸽇!��MEq�є�:�)��$a�3�&�O�3��	?�C�ozW>ʰ�C�v��J����n;3@2L�vw�j
����dl2_�t�y���Z����.�5��G<��M���B�G��g*��0^y��b6�)'� �V�
��� ��Mm�Z���&p�b�^+O5�~<��7 ~����O�pCo.f�~ǹ},�A���=|wr����o������V�Σܨf}I%�Տ؉}��$�Y���f��!��JӦ��K^3T��
�{�@
��T�:��ʊ�8}{p����.9cG���1�)�4�+��8uc'�J��HY|��#O��w�Y���\ �/���FYx5�5���Y�0���t�ƺ$fd/���}&k�5�Y8X�^��ˎRЦc��A���E�����Z��C  ڪ�z�	6�Eg0�e��Y�X��s%�sWr�Y�w��7F�+w���
^*��7�Oy��s#/L}:���p�(9;d #i}N��tva���ũYi���L�/�t~�ɕ&~]w�Gk��Җ7n:�s�?E���O~�g�gd�φ%~)��㾍�H�l.7q��G�Xx\es^`�|$����\�2ѽ�g��\�k����v�ݱΟ�A�:L1�������g�g:��c�����i�\������b�Fag��n	-�H�F�C-%��(�˃ h�T�>�J�������h�)�����&��s�h2d�P|eh|1�K���2����#�Z�Rn��
q� ���;�0��Ws��[�E#�=��*��������8��3��h?=����P�eb,ڡ��PSC-�y�a�U!|ɘKk|�;�����ھ2�9>�Ϗ��$�cј��\���k|�o'�-���MI�\�4'ȋ�.-�)_��V�e��7z�$].
I��eY����(?M��i\���P��:*����I�?~oy�X2�љZm��b��*rm[59�#S�xr)�bRل&j�M�'mޥ:���N��'���|	�����}5#���SP�Y����}x7!x��g��Չ���8|S�1Zޖ��K#�ҭ}�G,F��������:�jk�A�jf����Ru98C��]�	�[n|-IQ�{�2�X�ѫL8ݮA!E��e�#q.df�!�KŨ+�����V�z}e�f��&�}Ū�c��h��>A#8�4 �/b+����[�����#>9�ӟF>3�y��b��U1�:C3H��)�̰ �ÃQs�;�u�X�����>2�؊L;_)}��>��hQY���e|-tv�"4Ls���Z����{U��Lܢ|� / ��;�����\����/�mn"�ȆF��o��jB�-$@�� Ìπ[)^L��ނ2��׉$�d�M�VO�^9��w�K��K���T���N/�AiS�vv6�ۆ��~�"{1=�����yWk�����j|u����{�H�TGm�6w�mO"0�ߒ�+U"�7�G�V�y�.r�$Kb�\7&�oԏn�/�HF�����@dg�#���I��J��o�jˑ��gg�LȖM�H�aA^QUG�T,�``�:e��K\�)���ӅL]3�lU#�؀�l��4���q��ť����������[�Ԝ��������i�'�x����i�?L&��&8�3�c.�|cd������2���۔�T��`v�R
�i�vh�� .e�E*L�t
.4։�5��e�@�$������q\�|�)9�����}\>V�ښ\S˜�jց�#��\�WL�?��"O��ԣZ��hD����h� Yw�}r�z}z�&�F�TCj���l�4�1'ۖ"�E�$�:��I&*:����J����IH��5�W�zнut�e�����$jQd.�(f�=V��jAc���Q:�]������^���UV�b7Sq�0z��Q#���IU��ʜ-�{��o`��c�8J��\�b�M��]���f��O^C
 S���ޏ�%�)!K;C@�˜!#y����O��V!��n'����S������0?B�p-�ȩ �Y6G�8��uv��H���u��ok��k@�� )`n�Xi�,B��&Jv�3�� Ptj�H~ֹ���i����=3+&{��ޟ����03h�l-o�6�ĭT��t1A5�2�t�_Gu�pD��q�>�}��J�x�|���^��T��@�#T3��Î��^JT(�T4$�������B�_a�G�"��}��B�CO8�(�<ow��c���w����� I4�L}5�/3�70'UѼ���n���pl�,�?�O�Ȩ�g�O��`
�_Ph�����ԡ���W�])Eܙf��l���l�/xl1(�ͫ_6'�4!��h�)��`�*�fػa��R�:�V����I�^;��œ����n��+ތV �QQh�b��pi�+$���vV-8[<<�$u����Ǳw�j��ǋc$B#"N!�%נ쳪���^��z�U3�G�c.l$���&�߂W����|h(k܀�:�h�G�ɹ��G{��lg���}&x���q���H
{��#~k�A0	k2߸���,wޓ�;�+i�>0ä%��WE'
=dÜ� S���[��ڑ<�폳�����غ���O��¯���[M�vO�qsW'�G}d�Ѽ̰�0�|7i�Y���zc�����v%�����ˈ$�����7c��±��o��s��s
����ȯz�H�ɂ�{���oF�8d6��wA�-V�V�B	��F?�ϺՉ$ ]}���
�	
�z�v��l��;�{=�Llp�Ƹ�?Y�<��z:m�����>��ʔ�����J�[t�{|g�����(p�.a$T��k���Y�w�����L#�<�@�Ć��G`N4;���hH�1"V�ט���D�F��W+G�Le�H�X]� ���!Ge#��9Ob�ض�`]�oRԤ{�E`^�C��"���ѺP����K�_���m%iZ:��P~�c|���0%A�X|��D�]���N{�6[�ɒ�97[4U�#�3��-M�llT��>r �h��8����^�8��
!��<L� V���[~���7Oq����r�ƞ ��؞��Y�;K�~�;����~: j2R_#i��|����!ȿ���� ���3Dʄ]~��oyJ���"�U���\��Rl��Cj���)���0nHkG�V��V��yQ�������� ����:�6��mxSY�|����=8S=��w��YY�����^��tV*I�:Y����3v['�8�cUxpԔz3�O���q_,�[E���L^FG����w2n��d�CW��On���7s=�C<���C�
�I��8.�B�c4N�9l���xf��"��Z�hxl�C3���k��D#�Bl���U(�n͌��bٖ?�Ը2ϭ��L�T�q�,��V�ҳ�)�ϓq�g��s�Щ���7��]��F�蕯���Ÿo����8��ơ�����(C4�Wݎ������ǔ��Z7�p֟X��o�"H���I-�������#���s����7�V+
9�vRه�EW�eщ���aWO7�LI�l;�~lɺ��.�˂Kj�Q��;��B���|Њ�G;8q��ף�s�F���8V��-T�=?�%�S�oW��uEt�� ����T���{�ٴO�������֒��*K��Ro��kW�`ބY�I��MY�S�Fas��3s:JN�>�#���KZF�&,�x�䏾J�?%�ZP�o��}|�ҍ�bUϊ/S�I�0Wi���%�Q��g�?y˷�ק�~"2��Z9�o�x0Y	~.4�Bs�*���4xRWpz�]{�������v�^�ǧ����__6�g�_'�>�`�����!T��U�	)��9����W��r�r�{�����vv��U9�Z^�⬸7���O����6J�^�݅�G4���%���yI����yS��&{���z��֒H��Q��P���=Н%ÍS�h�p!뒢�9�Dޣ�1�� ��^�GGw�M@BN�}P��m�V��A�_���Â{�`��0�PNxy�#e|u�����݋�������n���D!'v^py�.���Q����\��<[O�XBVܶc����E�5��QoW7��;�%�����k���Rk�.��� G���0��[���IG�I��4��43�4����1I��̩�t0�%��,��/�z@8p�"����,�7��R��j��k�)w�I���//X�� �9��{���Jn�%��̻L�I�5�*����*N���ttC�ˊ�	U���I��4cc��LU��Ӎ�^/߉e��6�mN���}���0s���畡�^���S�2��iH���������9�#�p�g�H�� 	WQ�-�?q:��H?5����{tƇ�7��l\-ՄX�I����h�nP+l��w���_"�ͼ6�9(O��*W_�F�3h�N�O{����BFtk���gDU�V�i�vi�J��n�o��K�[��v�B{��>w���bU'�l��u��]��)�����x�)�M����~�k�H@%�Ր~��1~$�ҳ�Wb���Hȉpmμ'��G����AA�r����MD�Ɵ��X��Sww��Χ0
���Y���rY,�o��5�Sx�R�O����8���<�qb���E[�lw��?� N��x K�_�HOD�+An���r�\�-����`?Z�r�7zM� ll��I\�Sf�����Q�C��NjZ9��=���gwd�j,��:�U �Pdk �ɩ&'�?J�Գӡi���	`c�<��P��v7�䴷<F��T�n� �Y�v_ir&���@K?������V�&v>nu!��0�q�C�؛� �O�y���M7�Y�BN����\��ٵ�,�n��	��q��Yj%.���=�{k:��;�`��\�=�MS�P��?����1�8�Y�^A�ibi?[x�M.{:�PL�見p:��#��ٗ�.�Ry O@���]y�X�x�R;+�~�(�,�Bj}�q�jZCu����dͮ�<���-m�k6J�Ӱ�X�u6#a�
�`(@F�d�U���V#ܩ����":M�:�j`�����ı�C�t2�J��@�C���h������Ȧm������i���t4�u���Yk�3d���3J7h�7tg�@e��<�|���EN0�E����OBO�+=��N�����V��w��0��}�*��J�pϧ[?~T��Dum ^>E-�@��P]�������>��x�Sr�������m��s)s�Uc��l���Y{)Y�7+z�?XN�촺�q�Q�J��z+�Q���/`d���զ1Q����v!�c��Ĥ�U�O<��Ds/��%ً��KS�23��5�y\�b~���j5�j�hy����s�>�<MG��sf���)�Ϟ�V����E}2��oO���7'�q#H���qqW���;Ԋ�6�]GC� �lx{{q�HLҘ^�������bG�z�G+D3�͇��h��*�BʚS\�L�5�c����@J=A�&�Ò|�2d�30'C`�VS(�Sq���l�4Ew�y��t �K�̘y��Pg�2H_�Gu�>\ΐ9c��^�2"�2�<��SY!�����	KاB�������e��TLH�i�_����5[D��k�/m��)t����Gب0/��~qƙ�u�	|Ϫ��F��4|/�D#T8A@F@׻�e�z�O�͸@��?�37+�\�:��?�s�h���'��3K�<�pL�A�uO�����NH��́ޠf��׊4��<C�l2�;K��?I�Y���q@i�,cL-x�0\Ɵ��,��6�cΔj��a�o��=0��	�Sh�S4T���[y1�k$�^QF�9 j�E��SV ����֙�ﹶ΄lZ�(��ʿ]X���1��,8�HPrO���_�7<�������V~l!�l<b&Yq �V.c[�〟�M�9���c��V�^7��7d�1�'=��/����QH�����S�)�<��uZ�YBUߣkٲL��� 1��g��r$�{�w"d,�����|�e.��~/�z��Sߦ�[�4�&�&5*�{����q���y3�΄U� (1-6ϴS:���tt���wt23xUQ3B8>)�%�.���6�6Υ�rЍ�� �Aam����胰��pnL�;�S�� �1c�9W���7��F�S�d��߷A�p��L��
��	�V��^d�w���؎ȟ{�"8���q���S���Uk�.֣u��0�˯���q~��a��H�V:���Mf'���B����ˁ/��l��[c">F���(��;���8y��ڮK��d��\hI2�K�M�^����-)�a{}�`�Ѱ��E��3�'����}v�4������^Mj�n���}~�j}��7�ހ��GS��{`ɬ?#�ʷ�_��� `�N��l���._O۵?:5Ŝ00�M��Rj+���)����>��{�Z� m�JJ�����
G�x

��p�5�������f�A���c���@u��	U�9q�G����l��J�.�p�M.P���6|��RөV�ՐwG���s�k��SMS��{2F�؞����׀ӿt���-hU9fT�4.��iM`U��f�H�_��xXya��x"Ϳ��HėGD=(�Ry���
��r?Ըrg�*�$��W~�?r䑐y7��y�}�pR'�/]� nk?Q3�;A��܈S�,�S��\�#0Ȏ��D	�L�áhٯw�R%�F�ec%���m�I\����![�9����"��̴. ��Uo���\��S��awB[13t�"�:��a�Nxa����&�Il���Bc%j}�M�<�R�(G����e�O	k��B��]*� �y`^'���__��a�eu�"NZd��s�g#��os�W�����l�������˓wY!͟�>PXF����I�Cv�D��O}^����ȯM�켅z���p��O�"2쏋IX"	��xiq/��Z��9k�hTl׻9❕ݧ >�7m��`,���#֝�w^�I��b�B�/7����q�,�z��U�U�s��]����</��:p2_�h�����)���˓n�z�g�P[A�0ۜ�j�&/��坽 E�����e:��%U��"��:Q����,�lB�L� J��[�6�lI��͋<	/�������o����;��׷��F��B�i���9C���v?�:)���Q�z�0�G}q}m_��WB��v�e�c�(��ޅ�[DFEC`�;��J�d���[�i!��]������|A�2Ua� ]�@�!_+�� 1�v�ե�HJ��V����w�s��I߶��\j,Ջ�٪��u2ԑ��D��$/�s������6$x�D&{/����G��;.)\p�giZ��o���e����$���O�>�2s
r�=�+�^q��ƪ�kcj��v� w���oL�({�J�d d��W�gD�9I��?��;���7콪�uB���9d�uwD��H�
��.%2�D�g����=���qٕ�_�?>�~���5�������^����O?�y!
�Bb�2�&Z��$�{	9��{>���Y�41$Ǘ��j6�z�j�6L
{��v�D0�� �؟��ꐦ�F��y8��W]@��VǠ*Qp0�,F5����a��ZlY!V�O�u��D�
���`�xV+�i��<��pۭ�T����a�
�0jq�f��R�Q�
��D�t�.7�}�{5�WP���o�'�B�/�2u������2j6�q�2d��&����P�?���T�����s��~���d�M}O���rz�'߰��D���ڹ;l�p�ҨN���tq�ԑ���,Y]�(�v�.r�	5��\Yzg91�AZ�,��m9���5�>�4�h*�[���ڔi�:�ې��U5��Z��T�c ޠ}|�h��B�&aL?봮�� o���*��>v¡X������GU�kM��G۟�vQm���c%�m��v<͢�7�ϋ<�J���Izpww��k{����aűG����R��.���	UFԬ���I{���q���P#Ŏk�Cq�~���N�n2�Oݟ��4rȮ�m�+gW���ƶS�[��������|�	�֤��9���c�_ }N�^�w �Uu2vP_���0P|�xǫ\�9٣��.��j�qT򅫼�iG�gբVɘK�9�H�u�vx8D�V�q�$��N�Qs�Vk�ɑ�����?H/����H�p��R݆�i-U�7rr��v]��I<�/ʥ �K{R׾�>p������@�I��=?(���d�I��c4�����H0�å���=�����ףn��:P�
�z+,���Б�Ed�-�����\��t�|>�SHz�����Ѝ#L�w�I%��"N�i���OU�b�Lt_l�W��9Uܕ�
#�w�ᔬb,J���
���=��D�\�#\��!4���p�2w��)#>�����i��J�q��g� XF� yN]����F�Z;)׼
����wt�h����Ͼ:�P�H�}�YeF!�֎T�A�ɏ�r#M���|_�|_�v$�n�R�ר�����(��]*`��=�U7e�*���¼Z��=ۢ�i��g��ː�Z�3E���N+��7�O�eO݉_�0e��=%v���7��N�H7���%<�iz�7fj��	=��e�r�[:�;dE���aI���>���˒$Ó���'��xbeGT��};i۾���d<3��G�M��[����[B���M�`t�U�6�>}V�y�`�����һ���=kK�������vg�g?��r�3C�ܗ�DF~��D�}M��p��8�A�lM伞��u]�x��7'��*"���X�=ܪ���R�Z����v�*���$�m�1�k����*+��HO�@]�E�;���	�ff. y�����SF�^;���MR�S�F���s��H����0�k����[�o@ ����	�{pv�%A�y�h[��[�!ե�Qs�"��Q�T���<1�j8�K���<�4�r��:"��6e���,bh�*��,_-��f�xN�}GZ&}��I� -�7p��f� �k�w�q#/�X�F�����FH�EJĖl�>h4��0^_�1�*�6���e��qN�|ya���2�}�x�O���1BO�C�g�O-������_3t�\L�uIYiJS��;������C^Y�#����op��+�~��cæ��w�Kd'�Vab  |�2��4a�|`Φ]�O ��)#��ޗ,���*����  �<�'}�"�� �[z�+05j��*I*Ǣf�X�qaGs#��Y����31i+�+HW�OE.�����c��t�s��ɪz��
���(0���L{���)<��Z��5H;tTV��-QQ�m��'����̨$q��K���籀/�?����.9_[F�C�N-냠d���.{s�0dJxYھ0l�k�x�W��z���E��t2�����m |�6N�
�%r;��õ�	Z�L�U-0�xgg �;���YgV�0.�t�*��(��+F�;�\x�`;�O��SȒ�v�OC��X�YNrU�V�p*n]�����wVw��������ͷ'wO?�wN�������١)3�D�y��Y~J�J0p�w���Q�7�oN//��u6P>%����b�:�e)Az�n���*�����m��Ӝ�5��(�a �\�`ɦ���hk/�SdhYג���A��	}�&�#F?ǧ{��wfy.�P����G��8dق�����m�����K�,zx(�|�JlfOPT�C2�W�~67�	mE��V<a������ꫀzN���:c�{�f�Q8�ń<��Z�Qd���X'�Z��'J����Ճ��U���g�~�x��l�@x���� `��Ξ�w��B�&�]F�#$���O�Y��AE����c�p����w^1��"�f�
��b2�"ge|�C��1�~������kՙ��`��e�����
 ��h���8n�Xt�RGX(�I�%w�����ދ�!wlA_��ɛ�?&��`��´�O)u�c���w����3af,ġ�e�߇]��QCs�=5�ؘJ�zϾ�xU�Q��
�����K�#� G���j�p�H�#�-�#5��ϰi��U;-��O����
D�F�j'X��Na�m�����q�������s�b�&ĉ���X�DÎ �U�������j���".�Lg4�R�
vQ���%�4��i���{q��O;ԌC��T��׊T��iZk`ŨG��_WҐ�bJ��=}=��a� �!i3Y�0/W.��'D=/�1�[��^>K��a�^\�^�	����p����Cl�xN�L�LB�槔��Y⒥�7�ᕃ2Kj�/o�o�Ŕ*�}���~�	~e6����?nl�������o�c��Ѭ��c������aj��Q��_s��˨�I�?c���6r���������Ç̨�3�>Z�[�˹���#�"��E����$|O��bS%�w��k�P�K\�=�4����p�q�Y���;[(n]�I�*��z~���	�� ��f�fܗ��
(a���uM�T%;xI)(���A�6��8Ӊ�;6)nLu��Gu���=���!�`C��Eu� �pL��@�-�*��]�a�Ǖ%}K�3�S����Տ�Q��	?Ä�6�#��ȥAw<���᥀�z�tl��6��%��$7&�r��Z�����_�/� �9�ͩZ;G+���Q+��h���T ��b��:s��;��x��z�#3��N���	��
P�ⱍ�7�[/�6� v�	rG�C.F*�މ�ߞ�V��Y�H (�t���ˡ��ꔟJ�u5u<���b�[�{'>�
=�])��g�؝��	{N�7d�$l�#z��p����������k��n�􎶢8��
�>��&XC�wI�;C�D�@M|��s����t�C�W��C��������&��	�u���V���?D:v_�Ģ��8ϩ�Q"]�c,��V�
2͌r�yDc&�'���D�#�n��x����K,KУ��b�.-���6���=��([�D��nsI7�$6�G�d���y�C���� w�����yN/���X 9g�s�ĺ�9s��1��E�ךA�Z�a0˓c	 q�T�e]��b�Q��-.7̔�E.Չ#��2�?�<�}�j9`�H���Vڈ��n=����I� ��Km�-�=�v(�R|[�IO���݅�Mq-A����_�qF��%1���K�E�9 ׵$G��
6:�����FM�>�j;�.x }s��޷���qˠ��{m���w�7h��W���0s�^6��w|��D�!�E�ܧ��42����ߎ����ˈ��/����2d�������b1�M,���\eй�Dl���g��
��IG����1�3�5Wm���Q�����A�W��f�� �z:˄�-������R H �0�0y�8B���\���읬��W�A1?1��Ķ4��O����s]8�D s��z*!E��9&(�Z#;d�����7��ցI�o<�)���S^�"�ДLEs$�D�S�EeS	}�-~<�S�E32��T���|ɥ��&z-���.Ң�;����B
 �M�䭒@	�2|�E�X�2�����a��ק z"�(<"�J9��}���?�Z���.�H�.
~�٥��wlg��/>-R���`�O�Z�9,][�!5����L� !(�������-�������};cx�}ug�3'͹y�i��qe"�o��3x�U��B�G���EA�mg��fm_ǂ_C3���8�:�RxE'<6�c�������PG����?�2@7�VÁt�`�{������� >we�������������U�S�!<fb�!v�	������*9mި���?��P&�pw�����/�&3�*��l8=��`���/��UIf�l}^Uw�.$|ҙ�f|r�ܢ�^+k+I��+J�o�SJ�	�vs���;x�?R��˕�\��m[ �}�(S+ȧ'�/�t�!DM���J�l�\��X���@�$#0���f���Ɖ��8�Vn���Q3��t��V����{� �k;[�ox{z_�+������?�����ȵ����C�[���:HgW�gp^_zb~�Z���X7���J���������T#~�7j���LΚ��=��U��eW0�|��i�0aC<�#q�\/j%��6�;�b��Xl.?�riq$���TXLq��0u��'K\O\ah}���c�Th���C`r��d �Dn��N�W��
ޖ�?��}W�X�3����b�^���!x"�n=~���3�x����k���Ӂ ��׼��� �7���'���a� �֣�,��Xs�U�G���i����WW %��~}���^���*��#��R���d�
��}�'6۝ߝ����-�۩:�B�y<1�9��!h�s��v��������~���>����|�D@U��@V2�o`Lm�V�"E߁�e.[�>��%y����9�ѧ�b�H���<\�q��k)�^���E�_E^�yE�$��t���'�!�J�%K�p�/77D�PQ�7����*�<�� �p�Z� k���O�O��a���l���uV��,X34�~EM�1e���w��sA�L�AGɌ�� �w��W�{]�O�<g�aK��m�*8��T�H�f͒�
-�����5Ⱥ-IrK?�PDW�ƨ*���zbo<3��P�̾Mu^u����
���us�	"ӡJ�nd��@BR�#`.�	�%qbH�������1����w�5��	'ed�*'K��<�]�)֚��/.m"��%R_M\�$N�υ�,;�&E� �4A������Qv����A�ʲ�"WT�0�{�y�هb�'���\�!��G����\�7�+k��!���@
�0CMx��z6��L�u:�j;y�H���<��������H�7�9C<�h�筲-?�~oߛ��<���d�����E�_�5���V��X����@-x��Y���R�Z?Nw����ފq���\�wb��z�B��H�Ϊ@]��	���:V�l���e�,�w�V�����0�y�5�����1f���{o������L	,TT��|yWA f.��?ؒ(�X��4Ҝ�E4~�&�鍩�)��*'ı�3|fS�<!a�Fn������.�R����LvB�[@�%
�0(�xKٽ�w �)��{�L��.���T�`ޫ̸n.4@����?�����?�$;����ݮ�5��e�_Ax��ˁ�y����+�D��ԟ|���z����}ї��z�"U��?�q�2�7⎾˓�RX�&fA�x����$�����9�tZ�����8�SorLqH(/�/pa"��K���z���LƘl���v�<"��������|	�Z������ 	��|W��xRe�
	G��� x6��$Qԧ,�@��juS����р��)=F}��f����j-���B/@���-J ������=`��H�7"�327��5��%;�9�3!�4���11�>?E>�� ��Dv�{;4ӕ��GA�ѓ�MY	#���s �e�� �o�ְ���Y��i� ^SIݖ���+Ƙ��@�2��ѺB{�Q�C�g&�Kj�VY{��0��p�}�EޛO��B���
�C�����]��ATW+_��o��B���Ñ��\� O]��$����as��j��ddU��G�?��}!D���o���6~�}ob�S��� ����*��������]�M��|�u�
��v��f�;|��_<�V6����=��Z�>=��e�;k��� �7��ӗ�P�_�٠ݎ�jݿ��[�a�4:ZGǙ�{�Y3�~�'��=}��KdKZ|��yo���Ub�D���y���c��[�RbV<=���ڗ�q��$~;)|�<��k�#�'X.�g�����WFI��
���y���$�L�G���0B.y=�E�]oj�&`<(}�C���7l*f[����+'�EF	�E^�غݻ�1
-jw2�2�G���ײ�o̎Q�W?���ӈ��.<XX@h}��z�1��:fqa��7����/|N[��x���+��{+��Ӧ�H�p@*�d­(������]e�h�S=f|�'[����R̠M�T��ǯ��?\ؾ���/� (W���D���<ubb3w0���#��d|��Q�/�\kG�y\g=>��]
<e���б,w�M����?�l:Z�Y�ePl�}w�F3�,m�߁��@�ۈ�ri�S@��z�d|IF�fz�Ni��K��1��n�Ϯ���#bZ���D���Qޙ�+_d\��7�{�Hke���*��TL���-�ټ���pF�`��I3�$s͝�~p�W�2~J����F�ռW\M�h@U��_�U�j�r!��d��&b73�-1�½?ray����{T!w"I�//ï.[V�G��U$?= ��.��Iq�H*�������fY:?$h�I�N��Mwa��\Bܵ<�A�c4�ىy����gy��1Kzu�8m�g.����۫Vѫ����jˆ�K����<`C�j�Iu����J|�����u�U��\��8��Wۍo�������ω:/xZ�1^}Xu��G^���~K�W����awnS��xg{B��d�յ���pw�5�Yў��{����a��	V��π��dUYR�DH���Z'<ƃ�ޡ�8�̪/�1)�m:�N�OW���<*/�,�7��F�S��`K��͛G�J�/����\���٠S@F ^^�����^�s�p��C�#�"W���K|%FB�J@ik9#��4+q�G����pV�������0oz�79�)Ά�������4s�ev�P��o�>i�]�apǨ�`�w��=�R��DͮŻf��,;���|�ߦ�.�.Ľ�wZ8����Жjmc<7'!a����{m9w*�ձ�� �=�(�"�SqS�/T�$cs���7��lk�}�k�0�b�f]n�����K�ͬmNIb�M�Q�t�MZ��Zl42�5���W�c4|F�1����I��y��i�޲��J�ݞL��>ȱ�o��I)G�15��>C�J����z1.FME����*0Yb)������������vl���V��W!����4"M���CoW[�3NB�q�%O��W+a)�E�:v�![7���͜�!!i)��w�����\�WV�V�bO�){_8�6RM\���au*h|���$��kU�	�d��]���h�{��o�����u���@L���3���|��0������H��E֊�����-ҫdhFD��0��M��N7s���vT|�o�����W�~ja��.��jJ��'����c�����D65�_+<��_,^��w�A�c��8�s1��d��;���Np�V�9h�_��3�P��0t��<��'��im��H���K���|8K��=[��?���i�>�E���_Vy8h�I��_�8 ���2y�^���u��ȬJf�M�ŀ�]�;�?W!&��^1������[��|5:����X�t���[�_j���W��[�d���!g�ł-A�M dGv�o)�����-��Y��Y�G/� �z�g��wN7�)4�W�`�ן0��d5'�@X2����?�|2���dIZ�{K�?Ctť����xb">X0�gM�a��e�3�6����W��=��#v�=<�1s��ǠS���6rh$��	���k�@J�"�F���A�>[OZ%*(`Nt�W|6bA�ǋ
�#���Lx��@��-sϒ{f� $�J���jF����"��4p�R���c��psnT7 %c[�
�@y��Tf�j�q<� �6�X��,�(�y+�x�{�ߩ  ��K<�� o���(u8�g'әԮ6o�+���1�8ʧbޝ��6Q�_���B����0�`9-R�kp�!
����r��,KQTM�=BݹG:��-���� ��>��M��{�i�])�p����:K%��D;q�,�e�+`Sv����5C��H� ����k}p~mV���n��ί���?���T�%N{���!��D�w�k��
�Srnp�n[��e�0�����fG� {b�����mO�"ֈX#��0���I�����Ͽ��%o�ޣ
	f�"�ٝ�Z�y/>�G�j��SC0�Ӵ�(�,���!|o�`\�m���m�f�YC�|�G���e�\(Y�^3U8�y��,zƶc�`�p|�~z!�0�����0�x�W���u�����:*4h�,y�ә���a{>�-&9;�<���,�0v�3tbp�⛨]���d� �u_p畫����o�,铡B{nvY�R/�UW��l�
:Q�N�)��5��~�L�v�t�v����Q�	XJ����~��: 1
��X��[����c�Hy�+V�A�*���Rrϛ2v�{��Oo[�lv�V>q�����=��7��h�0��y�a����\r���nG����o�Խ֞c��󉊬�05sX�?���g����L��~r��ϗБvԱ������1�L�P��d0��Q���g�B�SM�t��8'�����*� �9���O�q=���s�@�i΋���L@&zW�c
�*�7�
F�A(��?��&�5>��q�d��&z���	*���w�*�B���*P�ZY5�.I�μ�=W�2����h(^\��I̔9̄Rխ�̲�IT~����;G��)Yi��5�!�l��}��})�
�\�ިR��x�P�ɲ.����I��3�8�GP�#�Jv4Q�YD\���D�ʖ���[z�y��Sr&�1��g:��닾,1 ���L�F��]`Rƒ�:�?�cl)#p=�_�'�a��ڪ���pw�����di	:����9Ik�aˬ��nq/hf��	� Y�����4�m*�K��f��i��߼`��|�u��?���￸�6��1�62�D��������muTr��D����ɱ��ۂ���e��#�F��t�V(�Pm�!��,�q�b���u=��VRߕ�k�78��v!�xQ�3�66>���˱yR��ˇ��T����ُ�2���& ��n�_/�L��:\t���u��Lw���(�$�k�����+A��O7�v�-�IA�SW�G��U_�jL�s�BK(��F���<����(�$�4�� �$�J�ߝ�Yb��Ϫ?V�� |�nh���,�W$�Z	�(����2�0x���g O+g�?��Pe��fs�^g�)X�ox4��s�-Q[Y�F_�-P�Z�&�6DRd�D�bc����Y����h���M���s�����yx\�eeqG�����F��3�ţ]O��7h��~�c��.��6[ L����Z����:cK+s!�r�H#s�r �s���3\��ܩ^�����ŪE��_3;����N��)1^	�bv�>d�AX���Rc�K�~n�G/����]���S#���b���� F-�J�����'BUvX{7[E�Z��Mx�cyjm4փGp4�����6�\�y#HTa���[s�!�D��N���|�����Ș���Mጺ����W/�����|ՀH��	�gN��֜��àp�}��)��{>�K#���~%�3 �g�5�	cE��m vSv��j��li*���7P��%`E�8T�OwFU�"O��� ȣ_q3�c\[	���g�ۥ�a��`_�zƥ6�|�*<�G&~��̪Yj՝} g6�w�%���t�B�H�(Q��ΖmjkÙ�lr��_�=�U�S>o�ϗó��	��v"V�Gi�gԟ���:�>_��	Y6!�!��L���H=�u�����2�@���F�{������5�Q���Z�����情��:�6�
�n&~р
,�i<A�`b9��+ծV;95��T�(�E��W�ʓ��cV�9�;k��e�������b��>n�K���P��n��cu.����aK��ޖ��:�_���+�
1$�u2Wz�]��F�
\mY�*m��ډHx̌�3: c�i/�q�J�����WD��+�R{���T�������tc���j�鰥l<�Eϑ&�o��{�c����<��V���h	���|ѝ�|���ۦ5�F;N*^K��m�U@O�6�*ۨR�yc�n��?��b�UK�u�b�����%�.���_�I+GLܛ5=����<S�C��
�:��|C,����5�z'fX��#��Z�蕋� ���IVʗ^{YW����C��88+�.J���:��~�V�6���<�zېr�_Ѷ9�p�ON�r��Ӣ�y���n�������� �^�\D��Wz���MɽU�֠!W̊������šL@c�>3��O-�N\�|�{�t�#���i����E �[<Pbf�3 x�[��L;3����g�����K���q�&��>
h�Yr�z��y�6r0�xL��i�޺4��ؓ����jҲ�̮&��f��vkL��1r�rx�����!��Y;Z���y����ӂ�$��������jw�O�|�[�jޜmV����u}��=}�}]��E��Ñ$n�ڡ���&��"o.6����:B�V�̙s��E{���E�Bz2]����BԖ!l�o ��{�u�RL�,�P��h�?���d��
/[�A���F�_Y/&Z�3q������N'X���a{�
�vS=����u�@~^�~(�T�,���o2��ю7臫��&�" �� .��B���|I(��=!T�]6�l�$���3x����ЮZWi<U�l�|�� C��;�p�w1��0����Fk󈈛}7�`�g���&j��ޏ	�Ԋ��o����Au���1<���n��G��j��
xn�����,��1�1D�3�V�M��?|6d?_3%:-1.�"?�1^a�{r�G�Ha铫�J�󤣿΂�����R���7��~`��#�n׎��@%;���6R�^��d���A�Ķ��.1�uݳg�vw� �F�x�@����Z��~׶����4\��~}�d@�a�O\g͒�$�T�a��:�Mv>g�L����Z����b�aQ'.��K=�:�6�]�����L;�m�k�E���G�+N͸�(S� �Ԥ\A���|���-j.쥦��X�G�
��e��o���f"��Y�w�ܼ�GIq�y2��}һuOhz��e��W�6�9�����/� L��".�i�
Af.��v���^�6��O9Ok�
]�i({�4� �'i�?Y<+;�3�o�JVo��'�������DE��G.ޟ����H�n�]n�]����m��?_�/��ٿ}�,��6�^ҡN���ڙf���67�N���,1�Sx2����C�27�g:4�����{�r2�]�^� ӌ��&H���Q���$�'�hd��aq�r�v�s�^ypbhtvm y���j(�8�ol�!P���+�X�8�~��1�]7x����t��Hr<�����<�&υГ9���jo�ݻfZO�HGS/H �K�+���N&���ς��[N�Z���d<�Mȝ.Ǔ���Q�H��^	,qz/q�}���EC��req�>ů�S1����o���J�(=e<��E}���m�;��#���]S_+u\I���IY���b������o�;]����ѧW���ay���w�{.(�u����1�L���W�����c}6�[�i�R��*��r��Ƞ�Oev���o�z^N(u5%tҷg®�����x	����S"WG=�͉ׄ�?8ʫq��DX�aā�1�|�{��,����0A����W�����RqR���!�V��Y(8=�3��g�dZ�@��K���ҙo�L�Q`����,α���ш7���HUd%$w,&�|�}N S)\L@�_��x���h��l C*[�j'���(촣�����\�N����?+�_$����\LV;Y��m�W��n�=���o}�U���k�YP��0=)���G������ӂ*��R0��	H�zL'A��N9�ڍ�I�1��4�(@%|/p�%~=6w�^�/�������}���l���{����I]���������j��L��q�ݩ,��6��~���l�`q@�{	�A��/�\<�E2�3:�#�]k7���&���� ^ٲ	;���p��ɀ�,dz�o݄����	 ���i�����6A�3����oo }�gG�H�W�Ӛӝ�Bb,�et��t��P����v eZ湔Ԫ�Iq�/��;�� _�h��:�!ǒ²18 y�$����������s$�ig��|����#��s2$㔦��B�*�����V9�Y�4�X�n ;)N��8Υ���93@B�$�C�@h@D����^���&�!����2v����R݅��ye��CUK�@�n�n �"\"��f�����FN��\M��kĉ�E�&X�B�-1):����ˉ<,�v��%��/V�@N��1�@��� $��C�e��?�>|�J�9p<)|[02;.=�� U�)(���]{���`#����I%�n�`���<Y�B�H+K��D�z�ӹ`\�nY��닭tO�ۢ!,���h��)x���H�2�Z������ �'�HP�ڞ�r��tƤ��ɨ�R�y�P����D��8$�ov� �̙y���dv&�e$�Ǹ<O�!Nʭ������`W�g�>�mNr�"�L�����`zr:��C(��
�Ayŝ(i�!�0�=�˪1��kc,Ȇ0L�$�<e4�w�fy��l'k''�[���Dz �	E<jC@O1'��u�_㎿x����&�������(ݿ1�-{��o~���l��W�|G�N�h��2�iUR�������������UK��t�-���W�m#WNW��.zg�"��g��o��oL+���Va4.��@A �5\��A_�YO�~�ڽl��%��Weے� �������/�c4���(�������1�w�x��~��G�y�<�)��B(�r ���� � ���T�L��d`"�w��3�X6��'�����%��3���/0���A`����:���k�h���6A�Ǫ����y����S�jC�',�;<�������bF��H�H��G��p�Wv�?�6#j�&]���JxċNs_���p�c �B�X��n4�T�? T�!��#_����B��!1��!Me�>��|��e��tI�\�w/�E��Xrm���FCCU�F:����J��9㓉���MXq5��w�����PSkF	?�n�vs��R�@���D�}qY4ʑ���)�9N�>��oA�|x���,�G*��:���*����J��柰��Lh�Ґ�X�t�(�����1���ө�C�b,�v��]�Z�FO��ؑ�<�G�k���5ü|˕�x0U��S��p�:m�}o�,u�Z(�_ʧ�ͣ�#��6`x�&���%=.�V�_��H�I��⁛�L�c�R�JAǳ����d�:�u�!��P�O߼����S,�oG�`\Ei����*�g��G��Ҟ�OR��}l�	�x6�@Z������y����,��V���c��o��jr8-n��`N��B�3�Ѡ8+�;/]��5U�Q��������*�3�쁒�'�[�ú�ߎ#y� ^�zև�G'�l���Z*���{k�]\��\��*����B�D;(�&٦&�A��u�u|ͬ�q�A$u肝b	s�ߚA}��$g��2u���-@�=r� �%� �ʥjD���i\<4)w>�n�؊���f�� \�53o̳�>�e5/�����{s
�C��M�̮��r��8����7D����'��h ��52���ـӮǒJw�¸~�
��O�@g��_ӳ��t��W8�K�md��J�|�o�8�1�ǋ>���R��[��1R��K�A��+)��|o�"0-�#}h�(G)B��r�8�Y߁�+�9�I��2Y,���ܖ����Gh,a���Pĭz�x����"
��N�����᫅��յ5e����$]F�[u�e3�������7]
�F\�GQ/����@�C�9(���5���ˡχ��&b��yqE ��D�`��q�a)���z�YdNcQ�\9����:=�8i���?�	֬6� ���o��<~��42���bt�*�u�H`u(X=r�J��4�B����/�٣����k����Տ�6���!�|mC��:ʱ�:ދ]Z�)@��3��	N�L���\N|����\�y$�*2�~4�jPZ��?"�M՟,���~��o�]����p?��ˢS����%�	/��Ly�;������$4�����R �t��͌�����
E�n�S,?;&	%}ڰF�~}T���ete���<d�\��h���x�o9;��ł��s���G��VrP���]��n��Cs��6ó�E>(}��p8`�����o���ý�m����B����K���z����ԥ�ƲK�^҈�2��W��h�W:�r��#�z�Xmh���@ Ƹv������N�[���>�U�b�Ҵ%'���Ɛ���o�����yӎ���mq�D�=�7K�ᠹ& �8�u��c��V��'O�7t}+��4Cr���#J��p�r�F����9䘹K�4d4��g(=W*WU<�x�(-�"U�z���i�b�`��K@
���}kZ�y�}�*,}a���x��Ӳ ���y�!�֎ |�N��T;T�]�#��L��������O���+��$"b
x��R@#��$e�Tp���H�˘^٩�5�w*g�po��S����慢Q��%|��?�R�v�1�2��#cCд)jl|FU��
l-.�z�Ei�&�]@0���@�����/|=��GN,4�1��bm����Z�M`ͫ�咀�{�o�w'Px04��*���Vx���^�ˑj�(����s�VW��%���\Fy��f����tO��ݟU��Z[0ib��3�$�X�ޜH˳΃]���'A�+��>F��53���a�	q1 ?�6L�����W��Wu)8�d$��M@ �5������F�� ٭"Y{�'S:U��+�p]t�w	�	�Rߨ b�=�d?f�?�m�G`���\����+��
�������o�+Ɖ�ܠ�CJb+�����4��zCP�4o�p��N����jآY��XVs� ��Eg�����F�F	���6�ޘg��_���'ۡ{�]�~mk϶Ǟ��.�5�EVw�F���y�є�'l�"�#��Ҡ����������T�a�GB&@�Ω}�
W�-ֲ5_-���%�A�8�o��A�-�9�ߧr���fb2՘�<��.�$v��N@!)hT�ҏ�כx��9���C;ԜU[���U?el���xe;��B�d��q��@xd�����n��y����4��Wσo��a4Hה�O��5BG~`�{��o�0���zf^��y4$��B^�0/���:u'Hs�z ���z��@�0b�s�_J�-�!�<#pؚ��a�5-hN�=!FQ�w��Şvd�*s�v�seMy;�����k������)z��J���~s���iٵ���5��c5�q���`���l��P���$��?+J)������޶�����.���'f���~�y�,�����	��"��Eg���w3ֱgg�3D�k���c(�,��cK��dOh,�e�d���+!YF�-K��������y�{�����<�=�QA��2�{���O�Q�[�_��$�F����>j��hz�䔳t?��7�������e6�>f�b�<��u&�~����#��i�W��U���q˷{
��Ge����R��T�Q�]E��W�'�J��)��߯J��t���P3��#��oK�-N��S~o;7�	�P(��[p����ɽ�n��� -��8I����zY~=׼$��a�՝S��tf.cŪ�Z��mi��i&����?9��(%�f�*��]��G	�r��f2&�r���/��
V��E�F��Oj#pUo�֓/�dR[д�m��ag�R���Ax$Ƴ��c���*yv:��ya?9��mi@b�(v��ۥ�鑰��맱ߧ۴�rwe��c6�7[��ˈ!��E��݌4G���FE�.5��N*���mΏ\�}߲Mɺ=��d�� &c��	v��,0Efd�"Ky3�����c�x����m�Kh�I�j���͎�3!���S�~��<�|�?�<�	xZL{�u������!�7��;���>���uu����KSL���N<�I�&�!��޺��0hK�7_�cY�%�����O#w ��Y`w����ж"��n^	1>�ߙ��C���[��&"�
��x؋����}���3'��/�f@wؖz*�Kc� |��P- j�� L�hC)!�L)O��M%��2�h����?3�+;f�$�4��"��a���άb�� aAÍMz�������^��µ���,�ĤFw7w��/�s\ESH%��T��lg��>��3J����r<���]+���hdMZ��3K�<�X������ϧ/$N=-�����u�1o��ջW�^W{�Y[�'���Zn�=o�C	��E��;N��E�rxQ��a���U����f���}Y������V�����oT/���ƃ�j�*��đ��^��sf`h�z�.��!|��Z�,-�7E�T�O�xv'�wf��{�1>��x��s֏6�;����De&_��X���')I��8��1l�]U)�w�8�&鞃�\�r/#b������-����G���睬��[\.ӂW��&���baS�/��7�5bOn~��U��b�d�l\���}'���)�Wn�(|�9Ip��/���S~�����_���x��I�o��i����)���&��[�~}/ޯ@ܕ������[��\O�=	�;9��:��x�s��> ��P I�S�J���6e@CcL��LMV ��RPoj�h���z��9r�S4� 5m������࠯%s����W*�:q:��k`JI�1��8 �FV�O���l͌JяA�9J�p��9}ʟ@�֫.j/���5h�������΍�ג�t�m\Rw3���\��9_����My�C���L� �����^gD�w%��e�����������e��>�R��<�OO�1߈�6?K}|g�rj��)Kq�� �����L����>�)^>]�6jL�J�C#�h�C��V�I%z^�ց#������&����9���u(�&kz ��򈟎$�����]���5H�O�r��Y�Rr��^/×�����U��[]�q����V��Qך���NQ�<�����pz�,���V�(k��iX;���U�&��읗"]y��rX����u�)�5��mb�8��!o�0��3D�!Lc#�k����3'a$Xy%J��)'��
�q�~iԒ����?ڣ䈦4U�>�IfU8ə�Ae���X5�s���Gl�СH��!V4I���?]�X�yL���^�6��ɛ��1�ߥ�
��5��"�������ǆ����XZ�0���W�ݘ�dշZZ��x��Gn&4����`y��L�O)���&�[ak+z�N|��o���B�4�ڱ#�7�8��z�^~�|�����o���PL�L�>�N�j������Ż�Qv���w�����7����ߊi�g�-�Cէ�0]����T�G�w
�?�xL�a�-�;$�Q�0����l�k��on^���#�O���$=B������g�A_R�C>�/�/03v����(5e�HC]���ឲyU����Z�����z�B)7���؉WY�Ѥa���(0�����|ZH�5N\mq*���k0���w7kFR�ѱ5.V�|�x�`�o倩=��cA�Ô�?2]�D7LO�.� %:��'C�H�v��Z��p����x�~�.㉾�c�Z�x\qfu�[H^�;�RI�ʽ��P���t/�j���	�װ���͎!_�C�
�e�������k��=����	�w���Qb�^��� J\�Р������zOl�ot�b�|�M�bՖ)��E{jQ�m�Q����rڛA��J�x��I�^��T\�.N��$	��ۓx����k��1)��y��T��3�-�gW�*�ݡ�*�5���"?5�!SUl�S.H?Q7��칠Y���װ/q1"�;s^����H��T����(���c)u��>��.���J�3hJF{�W]���=l?}ik&K�1O��R�"��F����򋸇��.[j�f)���[.�
z@��y���w�����G�$�6G��Y04�C/��J�G4nx���7�f"� ��:�n�#
b�y"j�@f�(ޠ"q��m��c�PN��W���F��"�)��~U��6��_��ְ�=🁘9�M��;������d3�녱��=ZC�g}a���طnV�X��[;�s��bjdPk�odۻ�#~��O^�]|�7����h�a��l�x�Ys!G�*.2�uk	0ډG�7������8$�yӥ�)�mQ���FQ�L��%+ltL3�Kr����֥��Zf�a�q�"{/���6�$1�U�"(g�����m��GG�5��k�K��F��5m����T����aJ��=�=�x�W�X��Tl%��f�s�D���e����}�
��ja��qv��i'b8�ۿ�p%�
���qMso��q(f�om��G�tU�r��<�\����X��	��{5������J	�_55�)]I���tø��*��%��2�g"q^߯���vH�t8�dZ�T0ZOeR���7�ְ�հD1%���g��c��Ě��Ys�w�9�QiF{��.��X�y�Ua�����vB�(�
�()���JG/�$�?�S�gyoi^������Q��l��.���r�D�ݓ���ן��B�`hpK���DiEϙ�>�P�S�<@$~��d�z}1��M�Wݕ���M�QHA��O��E ��GfcM���/0��K�|G�x%����Tsy����UA/���������4*׍�aJ����b��x��o��=r��u鍛qܗa`��;c�I@;d�$CI�Q	9��y4�Hk��������6�;k幺�- ��	����<*̈́����$����1�d��C�j��7/��^�o\��7��,��9 ,���X��%�c��<� �A�_�l��N~�}��>�i��Ҿi�d����e����ǰ�V��ɼKN�J�N�y���~C=Z#[*�>D�}S�d�y�&��K�G#o��V�B�gLI�������5e�1
�;g��_D�֙�G����Dpw	�����c	�eK#-U�G��x�w�������p�E����àL?/�����7w���ik�����5��N�-�r�z������8��U��E>~Mc��$���o�̞R����@�h
b�Z��I�$�0y����}8~m��������Y��{_ڋ`~Y���r����uu?�<u̵T&kG�rg��߫ʵ҃?�*!(�5�c![�JkT��� (���t�,��'�Is���`����to1+ �P��?�N��S�*_9�0py:�FOs9p���z�Q��>Vp�H�f������)���ĉ���p�ZXv��jvq o㹰�۳��5���N�C��	OA��|%c�?��_����׬�X����;���Y����w0�R5�PZ�ܺb��0TՆ�A��Y��7�s4lH0���=fzd� F��]c4�3����>���U��b�wf�@U@�#c�c�_�,A����G��W�;q^����yᆝ�I�ȵJ>>����^>V����9�X��	p�>ʽ4�����	�u�I�כ0R��}�5&W��I���ԛ�oO>��4���ژ0Jw��EBǫFT��MK�0�az�FMKiF46��qB���>��_��	����;��?#f��S���j�i��K�s�Cΰ�zqN�1���d-�Y���*>�ǆ�T�|����mS�a���#W����oi�5''|�Qk��������k;�>l��m]Z���Pf�o��t�vI��Y�)���w'��h�x�X�$�&�����
1��p����;�6��v��V�%k��7+'��Ո�]յsȾ�0x�
E���Q.�eIϗǆ�����{M��T�j��jTN���S��@O��,�r%7~��~I��W�f�d@���C��q��@Z~�KkU����C���EZ�8��ɖ�[����Ւ��y��A;5`�]U�´�����Ţ�L��8_�H.��D�ڗ�<�Hz{r������¾i6�<Q:x������wz&Q�D��V+��Eb��
D�/�	ŏ����
`M"q�&��u��2^���7��E@W�/����K:�sv}��nB�&�4ԕN?�D��2�iM����+�L�1�Zݽ��B�O?������JKI�8K�x��H=�m���ySU���I�ũ�J$6�����,0/��S�o�#d5o�fU�W�?��S3�����k�M�t��9>�W1_�����X��7k���b��};*��^�j��4���9�����iN	։7=wߩ��qG�3���h��7D8>�W�%�oN�}�^-_R�JQEi�~7׸�.Js��Jz�g���]A��s�z�:��Y�P��N!�i1�h)*z<��3ʒ{�綽��\Uh6B�+���+�8�����P��&��/�W�@R��\e�;�!�8�pJ�^*�Eu��57���PI�ݐ� ����o�Ff>g���^�6<��j|���GpN�q�����ştw��׃�F��d�m�nY�8���+��y�R��m���0;�1|ф~�#CLg�.����ݵ�����q��n�����)�1�{��y���N���N�0<�&1bD�羉�荱t�tT�#&T�H�A�*�D)o>)b�&*���1�&G���&$�	- _ME��-�O(-[{�+��
��LA�ГӾd����X�@k���᏶
��k��[��?5�

���}�q�إ�2۝O�C�����W�dϦW��7}}��G])Y�+����K(�~�!(�N�p�A�u���w���~�l1���X����XFt�(×�4+X!6���a�2+�V��V����6Y��'|����G����+��~����Lv�^j�@ g���֯����Q��=���.�Q�{g4�����H��#<����Fr�, ,�!�G. �" �Sٸ�Z�}� 7�~�|��I��%�Ö�\
�<��q�Mk�Ln��'q�2�/��o�i��_/.�z��(��nF�1���h��Vl�Fb�@Cڻl}��8{�YH�q��k̔�&wјE�����$L���'���V�Q�Ӭ֟�Z�k2��,pY���^����F�d�?��>Q�0�Pb峕7��~��ꔬ��3@
��n��X�~�ʘ��~1�i@M+e%Ʋ�����SO4\+�_�j:�dI���hV�w���@xi)[8�F}��԰9�۰��ӡ�����z�/DzB3�.GP�h���;��kY¥�J6>;#�����5��n<�i�k}Xt{���V嘐A����5g'|���mؚm��]
�6z����������ڿ��ƞ�}�~)�������L�X1<��$ߍaK-G���ć
����x9x _��z��O�_��Z�!�N�u��
�	 y���R����q�X&�r�-w���QnQ��\V+H������T~��PHÂ�:�W��fG�}lGY�_���8&��M����?t0PL1��/�&�����τ������$���7���1����/T����b����	��t����U�`4u����{�T_�=D�}��4��c�b���ߞ��:Onp֯�V�z�Th�h2u�l�xy��eŸ[sA�59<��m�AQ��R�J�[?�}<��KPm��+��L�9�D�u����V��>-���E~���$y�k"��^o��1�Ul�4[-�u^�Ap��t�3~Q��V����w��� � ��Jf�K�$6�n�
F�Ӌ�|.���͋�o¤��Ǭ����-��g-ՁE�9�{_���� ����8�Z�壿�d�FY�#�O�1��r�}{A��F����R�&%����,u�l��Žg�t�,S�N�:�+�b�D�bV����1A\nD���Ⲭk�w���	c�F���w{�Q`�����27�Հ[G����39	�(T����5+JF=�>�V��x�p.�GЃl.��G�8�����kǯ�,�F�8z��uC<$���垕���Z�=-��`:���M���vK����m����/|[�����Z�O��n�?{����?g�������v���E����6;�4Ș>����p�������ge��������Ս����^�}[=��}f�J_+���������+���9a�o��&O�MЀ�"!wG�F�_8}��9���k*`���3=���ɠ���Q�jZ���E�T?���:Is":�"�M��\���i/����H�|&�����f���]ƭ��y����;m�p�]��+���Y଴�N�=(G�(7w���i��ny��	V��W����w̻�6�J�	�ٔ�ǸR��r錬1w$>�O.�8�Y0:���k	W��������J�b����!���P���2��W4Z����=X\��r��$�-ĆS��([gK�N{c�� �6~��4��q��5�T:��\����ݭ�=p̖	�qf�4��,F�<������"��Vlz��@�8�z���{S�,�}�'Q���~[��tP��[�E�=y�`���o�8�Ɠt�3��d��u8���GjO��s ��
	��Ű�9G�t���VD�ĝ̴(ἳ,����@�lm	�nL�������Ph�d����$�ńW:�=����g�W��܎~�����W���PM?�+4X��E#��[��;9{&J�
�T����� ��	��1gWhH�bJ�c�jX�0���S�D��#�$�k�e�!+�A�&r�?�vI��J�ќv��Ꮤ�}Sf��A�X𒙍�U*D���*gw�F�HOj)����6?��"�VV�>�2r��"Y�:}��c^k����!Ox���ύ��5��ali%*�G��U���=TK|RӺ]w�*K4Eؒ�'�a^'0�g1���y�����4�%�����7�j�⨪�F#�U�������� 10qD����%&��uD
2���)���>�Rƕ�h���v��r�������K�� ��zYGF�i꾭S�{o��4h��>��k	K&�ʮ�2�1��͚������ڱ�����c��&�l��󀙄���ytun5�vk�Gʹ����:̘=yN�^�Ӎ�$=V��6��>D�+�a��9��ߝ�,�u)m�n~����V�>��ޓc?3�{M�����0)1�3H��D����I%v읯�A���!���׳�����[���L��."�S#��a����qB���[�jM���u	�@�/�J
���1������h0kr� D�C�X�}�� $����b<��%�eOX��UC[�pV�S�\���㘴��%�ι��ȣ�7�U3���i^w;�l��aQO=uR����_�� �,%b�=H�������Λ⡉�.Ƨ�_�/����AR\��\���0���:=�J��A-Ꝭ����T���S�O�X����BF�/�<�L����"D��20f��!�'�����$�V�(�����=ѩ̥�d�W�w��f�|�|�[��u����/�zY�5�Z�2$t���4GD������C�sb��\>�o��w�������\<[�������u=�,�߷tp`��w��;�e��/*޼h��08T�����.Y>@�T�0���R���S�M䥶fLr'єpp�KȽ����l���v\�l�]�R�ǫj!����-�vȱ(�S�3t�ݝ�~Q=;��
N�s�VΎ�~��EOi���i� ��+�L�{&~(J�)��	gH�b�6�m9.�HBa�����O���vN�6�BX��U6�U�1(~A|�rL�y'S��u�F�;Qڐ��k�b?^iӌ��t{n�<x��"�{g����W\�^P��<}D~�s�m;|�y��1Å�K+ںªYk|>�#+��G:��é)�zٽ|��svmj�����g�Q�v��gwͺoT�u&>��L�S��\U���Ϛ����j���$�{���\��W1X���Z��!����B*Pf�@�!����O�����L��H��S�x6R��E]ٕc�e��]"\V����^gΎ�D�F"H% �9�Re�锑D:��@��s����uH��Z�(P�[�t��\J�aڡ�Y�T��;�B�Wz@�j�:���;^���ȩ$�"���μh�U
�;��Z����R�lϔg%>�i%%����K{��됲�%��i�ߖ��H�W�q6���je��(=~����aE�D�s]J�z�n��9g~��kf�C��l��z8�����,O��'����X�w�\��	�Ͼb> �s��A�QI��x��9.,Eҿ����*�����G$[1jo�v���Z)z&d�E� �1�P����J�2���oV�3x_Jӭ5�5#���n��ҹt��!�����H��a�WO�th�B�xL7�|��J��4�$m��?�w��d(�I^ ҏ}P$hg^>>L[�-?���k�:�Q�3�U���W�L��i�V� ���>P�;Xf6Xk�c�ݜ�!/�3�CL*�7�=�Ҍ(����X�k)ɶ�Я-��.���[���
��Zy�v�(�B�d�:�oS���E��9�-p$����G���O���Fȱ.�U�`��&�L0���w����/��x*-�.�.%�KP]IGB���MI��/S6R8�2j���4������?eg�������N'q�����n4ztm0;�n�5I�w��k�!��jm|Q�ť�ә�<*�&�ݐ�#Q��ӏ>��cL��q��#��FUÑ������M!a�J42˿�eLGW(X�{��`�1�\Tp�ܶVE�t6�%����5	�5U3���I���D���H(@eل]�҂k��J7+�0Ah 6Nc�	�f[�X���X�B[���X9z��*�a�Uf��1k�e6L,^��[���E=������^@���ՙ5�Rb$���/J��q��Z�N����U��h�W�L'11���U݃�۩��;��U�N&����Fc3L�(��eBtc$N�����}rH�؄z� >��� @�{��zhӉ�w�D� }�5�a!�L/ҧDZ}���S�?QQ�g�~v��0�'�����.��W��Y~/2
>\�<1w'���h�(CS������X�R4��Nb=Q%���c���S�SVSS2�med�I"�
�':�B�1/��v�C4B4�_�q/b�����-pMI��~rY��O,��w��}�Ӡ��X�f��<!j��H�����L����d%a��Su*)�����RÖ Gʊ�N�:����yh��	�:���#�ی����䦡�;��O��W��@�C�TC��T-�(�B����* x�x��(���ﳤ��n����S�1���4G��i�\��a�j3�N�[�e����=0��}'�F]~G�+5�&���
�-둠��BV�X�s�=i=����Z�ɏ���Q�k[Neա$���3�hs��ʵ�l�����ʓ>�צ��/�&�?��=M������8��+ϫc�U�"�C�k�xQd��C؛{���W|=��X\��|��seoty�a?��af�di��+0��G��M���c���'���.qL���� [�&q�i�7��B�DDz�e7��W{\����PFB��8D�g�_��S�Щ�ԧg������*��]�D��O�b�����8���D��ߺ���Ϻ�B���S���p����M�U$7.�u�R��ƙpvj�ʉ�BG�L�"���WG��#@�JV�!�n���mp>�	 ٵ(�o��X��l�ĉ���R��{�N#q�I{�l���Q³������� ��84]V]jC�������P�!r[�V�4������0��DXF\1r�F
���d�X��ʱL`�(8;��p(����:�ض�sƤ�F�	 ]~�&9��\��Y��02t=M��s7�\b�\fjpe�F�f����E&��g�����Mo�v��[���4�s8z�|ۄY�F;����]o)k���~fcVG���x 9q���(`��g5̈�IBqϊ$����
�K\��[f�p ��<�Bb��5h$�i����~������Щ%qp<�=ŜU����6ti�[>���d%�g�Wo?��T�HI،)�G�ӌ �J���ޑd1�n���<bE�>�
�܈
�8�6m�<���2΍�P��v/�~��oʜN$N�1�b�c���<�.�*�0���1V+fL�η���j����lw
����@
�b�e$�Jy�B[H�4��&m�+�.L��09���x�ͺ٥;����E>W�I4�������zO?\9X�X:�5��\�p����Đ�N�2{ҫ95Y��{�O^�}��3���6�dN;�������2��μ7��Y-_���(͑���e�������ڽ�T+�|jm?�D0a� ���La���q"jýG���I8��Z�,P����;q���ҹ!�R��ȒvX��c��B�������l�k5|�OQ7��9�=4V;)�q]ҙP��zg�@dk���ZziM�����n�agk�M�p%��0"�X��Oh��#<�	A�-�oⰮ���`�f� ��9Cv1"�w�Lp5{��wx��
�k�Z��UM ��)��uӤ�3�v1�J�a_�aU��Rl�a���1���� �}�_�7�Ϛλ����qJ�l����V|�2B�J
.{n�D�}G���Jw���	���ⵄ1�"M�b��q��v-����b�m��v�e8��qg����y>T`�I��mP�1T-�tB�oaP%rg��_�^N�ר��8��T)>E� cH�$����k��2_��>!@�����  �������%� �n��[l����O����Tυ�U^DҠ �/ �=!��p���6��	6Uc-�*��	�/ W�㱄�}q3Wc����hq�YD6�Tc5�u��CZ�'��.�_5[�l�i8l��!&E޸c��c�Yg��R:T�D��{��'���)�Bz�����{0��%[��}�O0V�$���UP�J��x5!��@�޾}L�:N�������'v�}�N���D��@����Z�\���tH��%��w5������F#/n��n�y\��h���%��<���L�4�y�� t:�>@�Oݿ�ۣm��iC�r�w�QZT�Ć0l�*λ����ש��g�]w����������Q����5�_���L@����Tz.���}T��d@C^]h"2��]���c ���K�wK{ ��pFÒA���$�����2��,B7�_3z�����
������Z!���:� "�7�c�������9�BY��U6uK�X:"�4�l񇌷hiS�f-��m�Mt%�R��n��{&�]c���6:x�w\->|�_q�H]�>�����e�+���h���6��xw/X��o'�Ts8�(�P�/׻b`��K;�L4��	�0&����t`+�u �{��?9bL�%g/����v�FdZ�#��%fLiŏ�:����f�wc��tY����`��Ց���l�l+��B�/���8'15
z��������i=��;?ݴ����1�h*�!�m0�.��_�j�6.�X�yT^�w_ZK[�b˨�39�_`�g"q_�w���`��8��u_C�����)E"��_[��se����۴eX%N�|�`��G�h�2��"��C�����'��'�S N ZOT$u.�۫�^^;\��2�COt�Ax+"M%P�6 �]qZ:�#��BnB����+G�0C Ec��;qK���&����o{� �4um%V��-�$^��t?m9�AҳϨ'�[�^o@p��`��j]_z��*����}��(�}�����[x�Ň��?bN��C���L؆�|uŠ�K��Z�|1D�HOw(���ĘEd's%�=F���b�2"r�niȯ*���L:�=��Lx�T�.T��ӷS�(�����c2�ӿ�j�Y��ײh���B-��\Ґq�K��î���X��"�M�8�mP�>������� �[�=��gE7��xc�[}yEyޡ��_��nm�P����<¶
]k
zp��_�=��Yؾ��P��!��2�u��ݐ���uM���#��+�����#\������.���]�\!N|.�E�y|8��fJ�<�"d��v� ��щ�J����t?�\"�*!�����kuÜVGM��7q0[ =P�ٴ;qtB]!g|�k }&[�5��v�r@��9M�5��:P��2�Q��r�M�l����Ty�l�!� ��8�;7;�u=Q��-F��?v�a:j��$7i��
Tp{�j�r伦���~�&FuN��Yz赚�=VPu���_93�V�K�۫��ou.XCZ9˶��ۙG�t�T�ӡJ3	��91ia�����]�4�a���|�t���X�@"{�YDf��\|#�!H4�`<�QI��,K?P�A�Qk��@W[3=�:cP��1�+re�7�� Y"b�{���U�kZX�MK B����F�:Cq����So���ltK�yǀ=��C�-a�K��A���2�CID�S"��@31Cg�q)H�����	��O��9�(�ɰ�_E+�#L���/�
_L��gc�Ψ�vs���BwN�h��=��D�mO�1x	�j��^M=="�CW7�C�+���m�EDU��u;�]SFm��ss���Fy��VğrG�=4H�D�x���f|֯/N�s0�3�Ѭ�����E��y�(I���Q�)s���[1�H����"M^	`�G��_��k�'d�F���2=ẻ�u��]��\�\���u�3?�,1����r-)�xsFH8�Ozx�������7]��D��B�fr����Ԑ��E�x��1�[:١ua�>Ϙ���6����ٮ&���Cn{��)a�3���Z��e���]F#i�7��`	�q4ب� �J�?*���7���F �g|��ZI�8t?�U���LX5�{�m���{�������2ډ,��_a��9���e�Zw�_io����Js�1��CV��Ue_QB����M������{�[�^�����b }!���Q%*�o�_�}���be���Q&������Z��s�������	��k��2�R��GEcסC�@�:d����vtP���T�#�e������ِzc����<[<l��d���˷���8��Ky��;z�co��.9)�(�=^�_b����,uF$p�k��A���a�']'�!��v�v��^��G���O�h�� �'�o���Z�
I�L+�4�#ɉ�`�<	�'�4���P|����T�CėQ!B��8UT1���8���P#�rS�6XRA���ϝ�W�ݛ�1�[e�p*���Ϝ�֮���~5VE#��m�$�i
#;�g�8�C����I����P�&c�X� �N������l��?���?_>Y��࢈}`&x9v=�N[P�i-���K,K�ٯ��*Qڂ�' J�+�9�r�Fb��"l��jPw*�$Q�YF��Tɯ���#���q���� w�.��OX�T2���{<�r��*)d��b����٘�<j&
%�:���ŷM�'(���΋������v�?B��N~���4g�=�j��|�!³u���w�Y��F��ω��|����o5�mNh}�L	�֍�`�ס�Kc�S����Ҫ�;
�����O}{����Q���r�l����#�_В�툏���N=�m�x�uH��x����p�^�[ ���A(�gu���ۨdΐ�����w����q�u��؍�|9KEh�u���$gp��癗��[[������#�x!��ZF��nj����������)��ѣ]�Y�R��у��)75Fs�j(K�}|�u����Ĉ$G.n����7ad����ʍx-Vl�^;��E�S�?�e�Q�����U�>�H:i�A;�o]QP�������ПeG�"{���M(Um��}��M��n��$�]ˬk���!�uB���M( g9��]��:8���!E��fﳔ����F�P�E�V(����S`�4��&���#˼�c>5'�-4~���.b�gy$C������Ttޓ���-���Ǡk�|K�	�-�@���R�;"��R���fJ��$HkB��ey8��66Z������ͣ�qL�pb�0H"Cu'�F��Ib��n��Xfj��٥ĵ��0R���J��KY��Љ�Ă�t�8�\�^��D��	֒��l����jR���>M���#�?S�y�pl���V�,��kg�� 4WE,�l�@�<
��(<W�I_�Qde.N$	�/�s���S.��聧]5	������ZC%�,���Y�<�i��Шi'#��PR|��0���CIh{�,o�����m��#'�#X^a�pؖyAsA��.�ZL2�v^�U��cp�>��C)S�雿�Z��	-?Oc[7��V�'���ٱ������d��a�>B�n�N��|��*���o��v��������>�:>jo����񿉪G�gw���"}�$��X۾�������w������x;A�ZtX����ɊIV@�4Z*�)�4�G�'�q,U+��mz�2�~D��H��ѵ��g-k �pwĴ�~3b�:�Ep;�k�Џ~�;�����_�҄��tJQ�C���;��K"�"ֆM��� �%C>��(	n0�Ig����
�����[����A�o8l~˔����.���P�`�˞*Hx@X�]������Ę[�%�6��/+�<Q�bh�p��+�Ź
n5z`A����uZ��ǡ��V�e�����@k)Z[�]��$��P����4�.����a��	�_��?�b pw��8(6�H�N �V��wTp!�;�u���)���x�`�st>����5�yw���	��U�#��G��'VozZ�8&��[���N%�/dBX*��xz0J�*S��'��*L1Q
�����,��*ը�����T�Dr�.mxya�������U,��*M�u�-�<���Q� v���Ak�	J���Jg<ߦ�ב�B�f�N{+Y%�s�C�4* ���W>D�R��ƽR�q-���$��aPd���=����'�.��V��2�Z<K���~_�z�Qd��Xz6`�$���w��y�£��-�/DVeuS���P�yE �
4�o��n$ZgQ�<�^]�r`Dj;fn�\�a��0m���-
*�'>jH�\n��> 91l�)��z��P�����m]�+��B&�����su#u��>�5N�_�z|_ە'�ͳ�ٿq�U�ŭ���)�+jUe�q&��˥����v��=zQ���<L�a|@��F_���c��cJ�eȟ�y�j�2^׌h-zG� �U���U����bn�d-��7t���m� `��i�\�!T����l˟�XkUɺb��㔼���� 6��7ڜ'���:�c}�̝�M,�+���|�8�o�����o�Z�+�Se=�K���2����>����+-��F%<��~�	J8����>��d�w/+���8�5� 8\0�A	x�;� D@��1N�<J���t�10�u �V��+W9�~P�^��> ��jH�Õ��[ϐ:8(������֦{m����R�2�Fd��Χ�q"���̀n9 �-���o`�^(��Q焑s@�<	5�J\��>��Tnt����ꅁ������0U��Ș�*��3 `�&��38�N��-����RR�Ԏ^��Vy�|�C�� A
� �~A` �R�]�7��Gd�;8W����k��Y8N8�	(!\n�jK�@��u�ۭ�2ƈ�U�A����38�4D;nF]�JP&O8w��"�e��(q�e�q]��)O}�Q9  5��:���3�2�~�

%D�A�׵���/B5��WFR,LF���㢫��1���m�Q�����+���PL��'`D�û� ��|�l��U�2��n���J�w�E�R��Џ�JJ����+��a��1�7 "�����S���HePG>N	��|����H�	 �w]����~�= �!1��:fkHt�Gfl������vD�1p��	6�$H�s��r���UGD]������n���c���ﰃz��,~���`O�.0m�b��#K����x�N���C�-�����e�P�2R-+%Ł���o�m���b�6��b9���U?����,]k�V���x��jË���?罄.o��E�mX�h����5�J��f
Щ<�w(�`Ʌ@���Ծ������<�e��b &.�M?ʄz�j���O�6P� �4B�A@ 8g��!�(�
���.M�>`<���+'}&Q_��-8�q(K��M������}N=}��=����6�!���@=]y E=�٩�¨G��P@�9�<�@� J���p�ч�L���3Py"� [`�d�a�6n8��P\���y�pG��C2�zF�j{��%"ڮ��?]�|��a��QF�[�٠~'�R% � "8 T�h(3\l���8!w��҇��t�2��gf�B~��؀���V��Hh@ Q���PE��T/c�Z �2����2�@U���pGj�����}��p�*�1�^gV�N�B���8�(,�@��R;���l ��/p�� ��B_�\����~�{��a?p �Ѹ���o�n6����8�#d؄Qr$�|�S& LY�փ.9N�l��1H�"� �9�%���#���P=��BU�u
!�jT��� �a��s	$E��\�q��͠��+QJ��^
�Ͻ���+�Ku�:��pՕ��ub(ҵ+�<PJi�VP��B)e\q��L�t42HW@(�n�"�u�<�'r਽�#��#�ל�C��뀚�䪈�T��H	�'i7� �L��@`PJD ��Uc}����8�#���U��*sT���ͮ�b.�G6f�f{��@I��G1js��ٞ�g��/����l��t�Z��������{��b�Z��7, %���+K��C %�Zzz��u�ZM{���7ک�R���Y��l�����lz�U�v�%�};x�6�i��B����Y����Jl"�dpQE��V^[T������%�Ζ@��0�䠏���sD��!�v���nw���x>��.8Τ ����o����y�@��!X �Э0Q?�
�F�E0Ã����A�>\�2����9\�6 3>���v���}��bA� �YA�������e� �w�+@�&��[��[ D"���~) ��[��0 �%�f�P�s��3arU �s��Z��y�jg%�=
�>%�9.<����� b�Wfվ0� 7��L�A��~�N�z�ܓRNP  "������G`��&�R[���A��T�p�8�12o� Ĥ�2�j_����Ý���V ��
�zum�*��-�X ��8��>��P1�C��� ��A�O"�?���(�ED��k�������b�3�)[�� L��0�-z�Mԡ�ɀ	�P0)�K��8ȠrB�[��+������
�+P?��O���R���8��Zʇ3s;��.�C(��.�R��C�\E'p�&]�P�+�=j�~?��fn;=�
��PmB	QUD4]�Ad]�Ρ��p��\*]���n���"$<W� �zJ��CbP,
� �b�3cN�p5Qs�^.� rw���}HQ�PHa$��$�P� �� �l't(]�t9Pb�>��䪸�|�>��,(�|_������OP)�&Hc��c��cz6/����ٛﵧ�����߲��;�d�^����zd������V�z��3O006A�(ٲ�R-C*����j[���զ��,�,�;߷:ih��6��AACF7����ҭ6�p��R��*C8%C9��q򁣨�Q5�2��d�&��]n�u�0�2��ȝ..\uz����>��uz7�ԡs��(?�jp��qusn��]�B�m��B)-�l|�"�[�&�����	| @�"hG,�1�q_��To�:���sX�i\ʂe�q���@����<#�����~ C�\��J ���r���jP4<w�?3oc��fH
Mߥ/��sQA��C�S;��G����7ᰞY��Vo�]j3���3�����q�����Se[d�;�=�`��D��%���`�0�`D�1�6TF�U�?����e�9��Pb6�&�;��� 
�b�^/��]^����`p�Q&�*0J��.2��� % & ��H���F��ۭ��ví�jJ)p	�b����.�G}?�<���,�*�zz�1�2��!xB��-�r!*.TF@ P &J�Qg?y���g��S}�n5�Aqq<���t>ۋAQeL��8�thq��'( )��Z���9 )������'��Z���#�� �*�O��L���X����k��СT��y�_����H:�2�|.JI���>��~�]�����:�J�~ ��O���|@)W�p�A��@�(�MP
��BhQu�P��)1��: J�~$�� �O���p��gte �$)'�;RN�-㐂���
.��ʠW����h:`�PH/�w�������7�1��f���q��n�<�����ڏ�g�ߴ�{_��#oZF�^K;& ��o����4��U�$D���&���b9�i���b��m���fmMV��f�ް��Ъ��uH�+��+�?���ޚ'�Q��	ەp��$0��^�p���8b�1�����q��p�:�zS�����@� �`��@)T0�����1\~���Y��&t�9u��2�m�,�E��^���C�u��<�ץM��~�����(:\vL�DDnI�!J�]q2���s��C;�*�ˎ� ���������k�1��"J��(:w��.�M��������?�|&�J�h�p�`���|��:�����t�`�U={^> ��H�ph ���D�#,��H�J:�I��K@]y���
�3 ���&���Z����D��OC`!��cD�ѧC��	e�k ��.��l\�|}/��U�U/@��.����?��T�5R�LZ��0�H���}�J�e���>`U�lA�}�~z�K�5Q: ���@���9� 
�9ΥwJ���
j/ǉ�F,��RBQ�;��E č�Pj��0��h�=�)P'!�PR�)t���b+W�PY�QJ�@X�PG��f{\9	^�>��a? 
�u�!�l%��T��N0��bd�E("��r����"�T�g��9����"� ��U��!�HD�Y�!ذ$9n9������I9%��X�<��Y���)�M��vw�)���D�=ס�*
�<y���i��`�e'�7H)�)�s� �q��9c��c��汓����܅G�+���5�%�YJ/��ߋU�@��%Pb��.�SbBջ��e��K�0Þ���������W��D��}Œ���X����;#���Ȋ������}`l^r�
%Zs]�uuu[}]���o��V��V�կ[ݺ�s�6_�-�ߣ�z�3z�����zH����Fe�0�`wn&�`��z��a�� ���(�.B�±0*�:P5q`G�O0[sண}U��J@���.y=�a�a�Seq�yʅc�L�����(�=@�:��T�%�## �D��~ 3�ߏ���y Z���tp��J�;b˼u�� fm���Μ���B��M�6lX����EUN�@��$��2`	@]4� 0 �v ���Io�oP��&�(���C-����NF�A�@�zd�Jȧ�tnp�P��%D�[8�%��Օ��(J�vwG��]Ϻ_�sף�4�n3>�@�p�霠�i�o�i����� �$x�zsW]�/��PO�g�r����FY�pT� N�*�����A��=��!�p �8WNc��c���Ly�A i��%=w@��B��Q��P��N�! !̣j u�d�pn�Q>ԃ�. �}~�R������8PB�}J�%��t!z��S=u��!r�@ bln:B��;r(�*�N\p̲ ��T���$������p��C)q�+%�Kt��w(2 �R��BRF��P�5 �%j�S/��R��>$�D��^��N�A)9���p۹�Nj��^F��]uJ��,:W������J(����p��c�&Z�]�2H��)����`�	�R�ʠ�)�Jm���$_֕�=vT[�)^�<�6����`/�Yj?_��^���X��K��cR^�~��
XI�1+w I!�HO���xK����k���)���TKI����:,/�����U���BP�Z����}�&Wl�Q�љ�L�w��Z���0Bz0	 &�����hG���ha�}L��b��o` �g`���K�iJ�Gu�4���e<Y0P=�B=���s=�p�6Q/� Q/�p> ��Γ��3Gp��D��:�q��~�h�1��s\��k�� ��0v� 	���^���ud�u�V�qB��重���(���:���y�G�
���D���C�������],6[��`���=[���1f_hQ���G�퐡�	p\s,] %���뚽z�M:�;ѧ�!c^��nWW[\q��(��������p�C ~Q��08��|PP()���d8�"�> �C� ����6� tj�TP=CsY�c���͙���{�I�c{��?����`�8}B|�g��!Q/n;�u�eD�ݺ7�jDu������ !����Σ>(�p|�6A�[�\A��~�uP�QJ��)�tn�,�@'�8�t��!���@�8���x?��\��A	q�6a�B��5�@�a!��:����}��!B����}�T�=hA��Q��+��
��X� B�\��c��`b�"��Zu ��K��jt]>_ڇ��.�ʙ�gT�k�o@��!�sW�Ty��r#�u�W��2x�T�	���v����ϕ����r�N�s�nqe�(s�O��U�ʄ��fKM�	 (�R�8 "%�0<t�����B`���;r�;/I�%BG�z�_~��	6	�.P�+tD��θ��^u���Ǜ,Vmܡ:_����߰����mv��g,��.K9��2���0~����¤�V* Ud�I�$
Hi����`	qq���f�V_[c'�b�����Z�m���Z��my���>�k���ox�FWl�����zF)���%AD��]z2�e)�����?� �.x�ёѥ\�
����f_�6d8��<�`�}��E[\0.��	S�sM ���Tƥ0��%h}?+.D҅P�X����/u��,tr,Phk� !K��P������9�m�2r(ː㲛���\����?�<�XI�a�|�����ͧ��AL�)�%(1��A�Dұ�:��)E�w<���@�ǋ �q=	W� 
ߡ�o��j�_P�#`j��%.<��Z�|Ze$P[Â[<+GЂ�ݑD頊PAC�zl	l \�{����� }R-*��(�~����'j���6��a�5P������/��!Z�
b�e|�A�7/q�D�u %>M�t�]��c� ('T��c�x xP9��.�B��t�iVy_�U���}H���w2�(+�F��+P[���'���� @\))�<PA��>$T��E_�b� D%�pٹPuPh�B��t�+#��1ԑס}>�H�\�>� �Z"�Z	��.:;��
� P(�0b��
�8�0C��A-9�{���JQB�&P
��+�5R���gJ��@�B���eD�7pB)�e��(C��� @\�Վp
 �s>��9 %p,�%�.;���J�w�},A�l J��Mx7�:� Tѥ�H!�8Ζ2l���nU]D�I	�Ǚ�A�cv��8p孶�`�/�i��o�����3�՛�[��g/��{�o����Ҏ�̣�H�n+�B*�?`�)��<3֪rNX]ar��)I���hIɉ���i��M���a�����L���`�yy��_X�c_���lp�6&�ĲS����2�>�� (ay3�s%pMy$�;�'�Ρ�{&�*�s� J�`� ��R��3&�幉�_�7t� (!���B����z�`p��@*�P�j,�8�X�L�0Ё��s�2��9��<�� ��%��@���N� >�!,��E����\ۅK�>$�������|,�����e�^��{��b� j�C��M0��C������@�%B`#���� J����}� ��"� �u]��E���Z�t����.�s����pp��w G�	����1E���GR	������~�������d@ۀ��u��q=w��C��êz�O%��PEC��6D�4p��,�\�0,����3+�F�rp��	\�n���B�s8��b�\9	(��P-��z�Pp��Z�q8�}H�j[K���CDq�������`���2����<�Pd��(�pJ�@)�����8J�2a�PH@��B	�1���Q}!0�P^^�(I)��t>�S�@G����(�	�}%R�`�+���o��k�».: ������=�@���l�H;���d�qˡ�PJ�%� �K��,�
 4�y��2b�P¥G�@I�u��
��l�)k���:�	j �!l�� α˥���u!�B&WJQ��T��kfY��o�X]'��vPe�^y�i�@��?�h�޻Ԟ��ؾ�t�%���%��m)��X��=�B��cEI��`�J��&/��S#_H��Ӓ,)#�Ҳ3���Ҏ9dU���Tk-Mu�XSa���p��%�˿Z��_��J%=lC�dX�J�,�hC�d���usƖn�~:�y�fi�K��g���	ќ`P;N�(�A8s 6����1�n��Ӈ�!<����B�*�� M:��l0��`�EH�0��(�+@����.P[��.�yT Eqy;��U��a;�u��A�XP��5v�����t ��T�w|F�E���=z6��γeY���P8��CI����"���!�r��{S+�{*�hPr��st��|k��J��1��
�-�
Z��!�D���������$��R ���c$8�v#4��B� �Nz:�*����v�p
@�҈ncFl�04{��3,�oK�E@&-e *�	���2@�|���C>��Kk?��P�)��L[�����p~�� �|�����H����v$����tN˭��E �]�@��F�5J��]��ލR]��-��/28V��m��PZ��q����Q]�:�Y���FVm��B���V~-�X�S����Aʰ�vݻ�ɲ�Ȥ,uN8	��o\�"��<XBy�Uا�PJ�'�{e��X�y�@�u��PB)�0� ���\D����S��*�P�J
�D
�w "�(�e�\A����f�Tw���AɂE����#�*#�Zr������OR}y��� �x<�N��	��CI B%����.� �+n�%I)��C���"�PK@Єv��CH��j*AmH��IJI[��v�#���������W�b/_y��r�l{n�2���%v�WOYơ}vb�v�8��rbX��ݖ��ϊRYI�ޱ�ꬶ ��R"_HK�R,.%��3S,%#�b��J���A@����*kj�����ֺ������푯y���r��+���b#+�����ucZ��<g�1С��#\unHŀcp� ` ���+�{���۸ꡏ���@ma�1�;k�iz}Y2�2�}*w �6��FYp�<
=\Y�C�HPg�w�q�	a@=�0�#������~��`A   ���"�F�2���
�\�O�{���y&>V�;U�>5n:���z�.]������ 0 H �m��<'\���KR{QJ�W��@���J�J���/�A-B����J\�,�Ԥ�P��k��:���������^PG@+��P�3&�[����p ��9'��p�>�)@�%�Ƹ#���,�C8(�#(a��*�	L;�9 �Z�\�� �� 
���*� H��e2ܪH�0H�� �Cn�K�y��p�t�@5R�5]�~(�l��<.6R�@�q�%ˈ@�n��V#�4ݤz�d�B)�k��B	Ҏ���6C���A ��P8�}�k�c�=�٤vU�N@�����J��Q�o�m��	���P��du�R�^��� �|쒔,���TO�T�Ű��-�֕��P>tߡ�s�2
�Qv@�>$����(�G%1;ˍ�cq=V{Jz�+�yy�>�r�H��D����5�R����1G�KN��13[ ���̀zb��\A'�ٕ�@��t�K@2�9�$㟮}�
��|:�:dR<i���o�>�GB=1���	(�R,����'
0�7H�\�|�eGȷ�:t�|�`�ݝ���W)/��(��L��h<�#V t��������b�}vH��q�{�;����7��������k'�n��};,7�$�̸��+uT�ẙ�h���.-%��u��q��`	�SVF�e
L]-�
�*�����Z�m��Ȳ�������Y��/Yۚ�ֽj�u/�a�Z:����ʍ?o̧�nsC��f5�SK�7���a��r�Z�EP�?��#SM.���;�+1���bo��.�N�K$_��0�A���}��th���������5
��.��X J/}.�.��u�:��Q��|��*�Ar�2C�F��S��Ĉ2Kr ��1m�S Q'�[�6h���=� G��"`v�����]ǹ_@� q[%Ҩ�	p���0�z� ��|@!5��[m��Q�|Ɔ��*�.�8�Tu������N���h<�p�:��T�k3c8�kW��F��^��8��1��C� }C��p�1��'`|<�[Pc�;)&X1��])	(>.I ��d �T;��oBF�Ko��2�����2c)f��M���@8('`�ZFCs���� ���+��ZB�!E�"P; �p}�2+J��X	P�^��P"~���Q������o�:�Ɂ��J�t��;����s�F��X�����E}���0}�6��8�9�foF������a_�-RA�
0Wύ�l��	l_di
�ؓ�׾]��.ȵ{~�U��]�M�P��աkt�Ŭ���yA�����u(#=+�R���>w-��U��S�gF�C��_����ݕ�6�2��.$�U����3-�\?�#�j�$+�C�6�[kt�2�/@
��Q�^�lȕ�J���RHUv����9�τ{/��j��w��˙�Ae%���<Xf�覹��_��Ub�	V�M�� e*���M��6KUb��|���t���I�,C�I�Re�s������71�V���f�T�M���t`��ԕ �&�B�� DJt�e�[�qGwX�5�������`L)4�X3�����n�u�bu|?�[�����o��f/�_.Zh���e�����o	�ߴԃ�� �$���,?�����Za�aR]A��R�����l))I� (��X]M�%&�ZCm��6V[cc�U5WZmc�u֖[OJ�e��ז���Y჏Y�懭w�C6�t�M�x�'F%X����"���7�=k��[m\�eX��ȼi��2�l'eć���1zf����q��Ԝ�6�tR�
c��(��1��`� K��(���<`t��T�Ԓ�z�&*n���+��N&��1>)(QϠ0�9�:9��6P�َQW9`
��됧.��z�<m�zRu�*{R�Pzd�t<�s�u�u�.��9�*��D	�>�a�U�ȣ�h3��`���P�1��Y3���u�.�ie:����X(ÏQ^琢^�G�y��Q{�_
!�ԯ�˃%Fנ���]j�0�^}�c�p�TM����c�*GP�D����i��" ��:&$監�g�>Tn��6 C�2�Ao�a�"�WjQ�4�7��{e��C�\q��<HAeP=��\9�V���CD��;tD	vJ�1�Q+m��R8N	�Z��m׹����x���C�"��)#�!e�$0�Ɉ�.�J��G�X�����K��u��q����l���s���
Z��YP 0��C i���b7�����ꮓZ���[V���z��y����s�U���(��0�m�7�T��[/ص�*�2��^m�:��:@
���aq>A�h<}o>.	�� g�?&d%�a��	R�z��Y��\�����KCHa���<����L�\�g�s�}R1�u	�%R��WI)]/ �ٗx�� W8��!���wREłT��'A�~*�	f%7Jm�J*KƸ@�(���QDWϴ<���,K@J���-Ou�j,k"�`�BA��F�B�й�z�e? �-E�����r�:��;N*(]pc�����v �Lx�?�4�3�B"ܡļuJ�7[��Q�5�(�����.K��.;!P��y�c�����"�p&���x�={���u��K��/W��=������st�%x�R���w�$����V�c��'�(���H��XmA�5��HiR�`g���X_-%Ԡ}�/ �XKS����J������+~�ik��ϭ��bm���_���[���핏��A'eH��m�g�.�^bT�/!H�hM��MȐ�����dp�t����0jJjZF��0�J`Q�czGUtϩ�[�J D�<)���m��x�G��̘�O� ��ҭ2�k����2Ⱥ��2 ��-����V��$�#C����"���,8�K@�iyd�q��0 �r�ɀ��zD!����g�t:��zL�ʾ=;�IBFї1��8)�Ƞ�v���2�gF��g���pM����Q�U7.N��^�1Plj��A�BD΍K�0�Mo�(�1}Ǹ��f2�A����f�(
f@��0@_���CJ�Y��T[����tj�g%ӥ�>z����i��0n���^���?��͂E���R��r�ke�e���-�Y�Hߧ�[__H��=�"�O��O	B D�?(���D��zeL�a�1ϫ,m	�1NIߧ`�=�� ��7(.��֪��J���N�U-�w���:G�Ո��#��* S�`�%P���$8��Z/�r5Ⱥ��P�I�UG��i���V��A�z�oL�TG��S-�4
-����5 F�i��8Gƾ�:���&A�V������$u^-�]�jS�ꪺ�����8׬�"*G*MϺFj��Q35���P�e�D�S3nF�[���y)�:A���9�{���Z5z��ꋪ�:2���H�:��e(0]#e�|�5�Y�]j�JW�:*Tw�Tmᵳ�9�*n]b�jG�����	8�o�!�/��+O/���bP�1F,-`�fi������ʸ�ndȻi���4�(9�dȃ���EW���, %�ÔB�RR��<�?�X|�>�`���,U�$M���n���0���L/��Y���Rd>&	�SI���?DPԈ���(^u�9Vu� >�F��L#tL�Ơ���S��ê��+o�__s���d���e�=��-�g=z.q߫�u|��
D9q]��XyV�UK���MG0�5�XkyV�))���t"���eYcC�uu4YIQ��=`Mu�(U�T�m]��H��Uv��Ѻ��ىo���|�[V��+ֺ�+6��q�Z�et~�C�&�)P�H����|��^asWɈ�>��\H2�c2�#�E� 2)>-p�d�Q]��p�a@1�A��
����z[��Z(�>Ooi3U��4�l���B��%����;�F)��!/s���1
�f��9�u|�O�΢M_
y �;L,�_���P�qg��t����EF����>%��P=(2T��VwW��=����f�.51�<3�덜�7��zR������l�'�7`�v�"o��\ݿ߯���^�
H��'s�$��5��V�>��� �)��'H�L9�hۀ�K3d�.�_o�+dP���D�!\b\@^  J�dH@:���� �#�>��AX R�Z�J#�;����"��EϨ^*�R���D�m�Ρ/��CRn(2�C���_��m`\hR[=r����Z�L�f|�6a��3xVu�'��̼�w/�)	7J)	���w"�(Ϊݡ�pk5�M�Yȳ�.̲���.�T�ڦzpW��R��e	Ե0�6�'�s�_"5RN_��W��T��7 .D�F ���W��r�
�{�^�t�-R��n5�h*Ϲ������U���~q���Z��V/$�W#�]��*�� K�����$���>Bș?�\��@	��p#V]��q�~cˬZ
��9�5 W��̷���j�%���+U��Y31j��T��X�v����
4Y�
��#_�/�Vq��˖
̼v��B)�|�{�~ijo��P�S��M��n˔�ʙ17�,UJ���Y7	z�N�>'K��Jyd�� ֙� ��.��y� $`$	��	&3�QP�󹎾 ����Q���̴ �}���bqR9(?.P�]E��햢|ҍ�fP@��i	7�tt\�uD9��,{B0#����~)��S��yH ��}��<�v��ӗ�h���v{v�2{j�R���ն��?������y�8�Ӳ��F �y�r�V@*ˌ�M�0j(J���l���-E)�D���YKs����K)UZ~��4�Ҿv����ت��M`�,��-�6�,�?����{V��w�����Ц����mr�vvك�rFelG������`������bc1o�zÿ[�p���b"�TF���].�#p-�� z�/�`C2�݂A�U6, �,Zo�s��e�fː/����λ�$c��O=�,�} kX@$T��nK�3�X�\��)%q�(0���<�9g�몾.�nLǁ,u���8�{�۝t�:�ƀ�w�<��
{(܈�fRj
��#谮�:����>@�My��`�\��z=�O��R��`�:�#�B��-xҶ~���|X�[�]R5j�lە��|)�%�1��37 >�Y�%<ߕ��J0	�}�jk0 7pҏE�A�q�u��d�GY%Vy@�7���,�1`���1ƈ@����WY��ˢ�f������~u�γ��!�G�^:\��z�ճ��[(+��R�2&(#���gJ��Ol��A��N�ʀ1N�Sm��q�����=b�!�D@�{dv�F��6�K�Z��j�U/+���Q��e�ۦ�O�~�7���~��*�&Zs����h��r�}:GmQM��Z������^J�� Ш{!5��� 4)_��aF�z�k��U��qI��;�S� Do�5z1i�o�}e2��[������\���y�O�@��8��OB�+�rV-�R�қ�*ϵ��d�Kex�o��T�V,C[}�|�S�ʛ�Y�x��f�W��%%��4A�S�s���`rU��d Ё��GR�uj�~;e��K��@Xv���/+.��)��)���(	b�����,��y��n\�2�*T� W��Y�5��������6E�����}���uo)�I�\/0��ħ �VK�Q
i����
@�`(3fY�͂�@�K�q��K��h8�D��T�c����'�&Tͭ{�8c�%�4�b����N\ό�J*�2�.�уPK8xD�>���Z���U��~Ǉ�?À�W�g���Ϝk�,[c?_�����Cv��i��vY��]���5�:��S^�>+N9�_���i�sT�oL�:��J"�BJKO������h5�e�����z+�ϴDA����zk*����j*�������;��gS�e���[�7�o����u<�oz�F�<d�+��V?$���e�&��?t�X�<�Y/Xj#����2��K��>��.d���
\���p�
Z,�h�uܫp)�aA�ԭ掻Jm���˷ڐ���\�7�Uvz���m�~��Y��	�_���q�)�nH ��fDF`Zy��2d���Ǣ�i�q��+�R��y��l�i�E�:>������
� �zBF���u�Fd��Q:2vȤ��OKЧ֥����O��l���}@�yZ�gJ���ا����
�[.�}3pt|�&�Ŭ��I��X]w�(�;����,K@	Z,����r{d$3p�
�����=d_/��PD������1\~�R��`�)G�"�:9Gm#J�F�SP��~"���n��uX_�MF��1=&�m��md(9�ߣ��ֹ֤�[����4���v�u�W�m��Y  �s˸��M�~�`�ɥ��~����$�n��X��K4X���,�ʴC2�D!�%�KB�RҮ��(cթ��6=�z�6�~�Ju2����w֣�V@j RzIpx�{(�,c�*iJ�n���"X4+ժ�Uz�mz�]���k�=W�5�{��Aj��G�Yj�s�8ެ�i��+��Ԇ�uG먐���3i�3��ث�Zu�٠�z������t���$}�Dµ��j����"��.Aj�`'@�t��X��&��Դ�S��[�X��)Qʕaϑq,�wX����ٖ�}zN���l�m��k�^���B�	-��:�R*L��ؤ*��
�l5��{���*U^e��")���`��r���2�|��2��P��w���X��{W�8Q�� �*)v��
�'��q�#/]�?��ۤ�fY��~����[.��B��r�/]j*Mp˔��O�����n�}��2��県뤦��T&I�A�����gF���;�|���YȫRK�jo���*%�tսv\��Q����3��U7�of�e���~�b�}o�����V�o��gI{^��c{���Y摝��x�C�Jӎ{�7@�̎�+ ��N*�RjZ�%%�YNV� Se�z7�8������I=a}Mծ��Z��V@�n����&kmj���&�η�Wߴ����g�{�ֺ��ֳ�a^���Z�[���d�ƥ4N/�dS˥l�қ�rG�W��,���g�-ձel`�@u�����x.�?H�Fe#�?*��oP��S2��dL�1�<%��vH��'e��d�N	(�:�}�W�a}���=�d��0K,�����ΡSY�T[ ��YR<ݤ�0��P�_G��4}Wz#��?���IIL�0	6�2 Ȕ 2,��/��߳�N0�z��c����ʃ6�f����d8�oB�`\i���~��}�T�]j�):vR���m@�%ݙE|�	Fe4���CXzd�X�pRy�Y"�qZ0#zLƖ�w�i���E&��ՀQ���Ô �u�AvT�e�'�H�Pv�!�� `�z0�@�gu����sB�w/JJ���v��L�X�3��O��0Ȑ=I�KףJ߆��1[��Q}�{� d"&	�g&y �K���T7�Bt�(���놳B0_^8^��{����9m���.\�f/�5}����A�	�Ƞf��[�v��]G9��$��CT'����8��.���H=��Q�&&1��O�Qy����n�f��1$�<�H�F#��[Y�i�ڥ�4���T�� ���꾪��dq�H����ݩ���¼~U�ܣ��kI�]7���ýJ�;�#52v�*פ�끖�t%Pճ��wP!����B/(�R��H��T�)��-x�e���B�+�"�)��rh��Py&2-����Q;ʯ�Gmo��ģ˕g�U�ML�$�u����ϥ�Ң�g	H�y�ʥ���Jd���,u�x(���(�f�	l �L��e�$^�̹>��d���|wy�E������/W�f��@��O�D�ǳT>K� ����W�f��|1���AJL���B�%^q��9jN�yҕ��B>[������v&���O�^�~'%��;�=�~�`��|�f���Z��CVr��F)�vZ�R����^ˋ�k'�[��T�y��Ҍp l���Jҭ6?��Ӭ�2'�Ĥ8K�B*-η��fR�@��\k��VQ�kIq���$�Zʬ���Zk�VejZ����ښ��F�lh���K�я,�kߴ�'�i�_��5l~�p�z�Ɨ>`c��T�^N��b�W0M3$� /���T�[*7�(n4�]�����[�d�e��q)�i�)�0���̈́޴Oˠ���_jB�O������<Jfz�&�AH  ��i�G�y� AjL��o��(/pVn�S(0�t H��}U��:��u6���.�3��z{�����&�de�X�|z�V7�tO
�>��דқ���ش@5 �&t|H��{��F��U�����3�Vw��7�ob���ʪ=���}�)��;W	����u��X[��XR���3�h�z�� ��g�3��Xch�v,��CTʉ�{\�zi|bW�#TP�'Ƙ4�`���t��^L�`9��>Cz8�pt��ls�������:�e�Yߑ����	J�L��V��Xb��f���+
g���;�3�uU�0`�~�Lwԣs1��#}G���1֔�ʘT��a��Ԥ<}[Cz������g�P�|�>1���d�Ttꥄ�L�����X�:7,��[���k�Qm��~����{6�eA�o��1K�A�C� ��_l@��.}O\�E�:�f��3C���n==/f� d�e/}y�6�&�t�E �R��T��ٙ5�Zj���v����4z8�
�{����D D��B� �:�b�@V�vU� V)5���J)�\��X��e2�5��빦�������[J}ϥ7��>)"���)���H]ζ�k�K�.�`��+��a���d9����^��\n`6��YGb,Sp�K�O��`�R��%��~��+L)��k���	�,Xz�\o�a�1ϝ`R��
���2H����9�
�`R؋	�V���R�	�`|p�`�2P" #U�	e����|��kYe���{-M�Lӽ��yY�ߎ�_�n�?���������s�ً��+��G���~������u+M<n�I�,��nKVJ�:�<��2��C�/ %���#��@RE���B���k-�
"��2��:W@J����DWG]RЇTgMRD�A"�;?;ْ�XuU�uv5XM}�5w4��I��-�$(�6�ڰ�M��˭����w�k9��7��
�<j�[��-OZߚGm��Ye�O�x@
�7�2ΛdﷷV<�o�m�sj�6�W����e����mXP�Y�٦V>d�U��M6��~)/)�U��l��RL˶yV0/��X�zȆ!��  A��T9z� �Emd���!(� &A�<����H�c+�A��A�4��[�2s�-C�ؠI�%Tƛȴ�e��"C�qir��%h`X��IPO���VM�˸�Ɉ�E_��L���UO�����0���Y�f��[�"����%P��vk;����C6,X�\�ͦ�?�z4����q�otɃz��[V'WɆվ^���g��ӯ-}�z�}�ˈ��v�v��6�腣�����r��֫��6=����@N�7���~}_��H��	�]|�˶�:2���H��s����1�Vz���]kmw����~]�v��w�EP�^����yf�����=:�D� �ǋ��S��g�T[����ө{mV�<�^�8���`Z���u��M����SϠ�Џ��[��Vo�wס<紫\�{����[om��E/,����C_M��b3�V���ѩz���y��{n��m��L�^@��n�VA����[�;k���8��v�[�"�Z��A�_��K�@G}2��"��<u�[�Z�:)4����y���A$��U�S�NP��B�|:�Vu6�լ2?�2��E`l�9��f�@T��-w��5Vx�v�-�tm�u���Y�35Q�@S�v��I��u��0�J`�նJ�����Ww�2չܪ�_���Y��Z�]��T����n�o�zi*�k���*�T�R��Y���Y���Z�R��Z�TX��e�/peI��'�X���	��K���O��`�!��@9ڟ-�d
R@قO���+��&�e��RgY�R>����(+p�x�@�9�/E�6�~,���*�͖�ːҌ�H�z�`s���z�'(�J�x�t��x�{�����;���s��s���.���.�oϽ����',g��V{�r�I��6က���r��\��<���ﷲ䣮�ʳbH> V "���(Y�(�þ[�3��&/����I�N���-p�56Tz_RsC�G��וZB�aKN=nm�u��Xe-RG�Qc���"�����Wk�mu6��dc���xp�e�����-�+߲���Xẇ�|��V�T���de�O
k�S�lg7?a�7}���>j���m|�c6��Kֳ�A�������^�ӷ�a�]�}�<��1��Z�%%}������[�����[����#���GʧO�X��2���.�k�zkW�6>j-+�X��ڵF ��%�^��u���}:�[�n)�>�9�z��h���/P�^���(C�ox��hۯ}�K�f�>bCjC���f��u�u�X��x���Z"H�5�͂c��ں�����V�&�Y/#Z+�	�zv�:^��[t�k�1l�m��k���^����X�I m^�՚uN��h�5괭Q��CϭE�ؤgQ# 4��-js��Q�6�
ʍ:�I@�W�k��,^g5��Z�>Wk[�d��.]ouK7�m2ԋd����5֠|�R��^���^���f�j���ʪ������
=��{���Z�b-,+��ZʵJ�Zmc[���R��[��ER�y2B�R΅�\ ��K��s��) U��%*_�����Y2nR��s>�H�3�Z�]20ڗu�"�Tʽg�e�Zbw-������R����U?�)���rt^���L�T~�m-�Ŗv�˔��T>Wj$K0Cj!G�4��.��)#�u�����P0k���|�K�8��tՑ����f[����Y��V��I�yi�,Ծ:>�V�-�t]%՝"����Y���=/×p�lߒg~37t7ζ��\���������1�����}{\��&ʐ�\���{-^8A�%^)Y�:]�5E�`*���
��ʬ�R%'��5��i�W����嬠* ��z�\K�Rm���W�n����I���9$����^cI��ݱ���>ߎ�\l�[̬E�2�%�Yn��]&�s̽K��=����Evb�
;�����m�-�퀠E����c�.���z������<v��o�ݯ_v��~��J��v)��R0{��z&l�|��� ���Y~��[�j���M�e�����}��[Uf�>�io��:�뚙^��W�n�ٯ��Uw�+ʿz��*����^ӳ�~��t��s�ۥg��,����w�-�μ������6��W������-��g-q�s�q�O�'�����e�M�k��,/f��&���=V�*!�gU�L� �$YCq�5��Ycq�uV�z?R[EV ���(����E��&)�f%\v�M5V_[j�͕VV�gGcu��tko����k����&TU� �`�]M���f-}-�=�nC��v�����w�����v��oY޿��~�_,o�cV��!�_��j�l��e�p�˝/�d�/�`e�6[��V�b�.�`�k�F��V�z�蜢�X�b��p�ʀ�,�d�2|��7Z�J���MV�B�e�d˖m��MV�T.CHb_�����WY��jʜ%�>Oe��ɗ�ӵ�k�:h��U"�J}�KtL?��yz�!.��-��Tk�
��u:�z���Y��k���>*T��V��+�[���Z��%��T�@�o���U�{-Q]\�D�.Z��T X�.Zo92��y>�,_��9�υ�6[�ߤ��[�d�V��f�run�>����U�[��m���J�}T���;)�s+D
�w=�2�Q"`�M�z�<��e�k��Ϫ�V��x��жd�f�X���m�.�l������o����uѤ�<L��͔����z��=`u���M[>�/�6>lE���U[�@/��&�V襦T/7�+P����>j_��m:����)O���s�sy�����x9ʗ��b���ǋ��R������\��[����s��o'g�6����e�^�uO���[ކ�o�e�Y�������9�?M���P����P�A�ճ�Ys���8)_�r�>`��������Ԇ4��2�sTo��m��{��e��9C�MQ���}ǩ:��Pu��y�������d}�I��HZ�֒�{OTJ�}�Uז�~���-�������o-^�b���AZk�z�9�k&��xmc,��������]���N����M�y'��r|�J��KK�<է��R�Ǥ�������� q�c��!���%n��Z����j��}ҳ<��;�txC4��3ݯ��ȆGm�^<��~ot����⠾�~=�}J����C/��ݷ�v.Pto�j�.�`�־�`�v�]��w��=�=�/�>���V���7f/�7�]f{ul���Qګ���짼�N��������Y�M�>_�􌂴���Wd[~3{����y���K��O<j��yʊX�����~�uK���z���yt�%�B ���
SXF�+H�'@��Xy�a�g%���X�ˏ��B&PM��Q�2t��ۮC`����3�}κΎ&kk8���C����e���Ӷ��
J2-&����Y{c�u66yjoj�:j���Fk쨷��fk�Z{Z�O���3�mv���Ʋ��h�u��o��>g�?���|��,��_��/Y�+����-��Z�׾f�����=����s�_��'������e}髖�U忪����J��/V��7-�QI�Ǿj9�>n9�<n��)��W.�쇾��e�~�K��mn�~��T6����G-i�Ö��,�/[f4�|Iu���Y�'}������T�ڥz�t�RfG׾R��R����5<�Mk�Z���-k��?[��W>���}�[V��oY�7�i�O<a�Je�����R�׾aeO|Ê���/�X��o(}ӊ��+�}�E�����m+б��|�B�U*x⛖�ķ<�_e
ynO�����*�h���:u�j{�W�����k}�JH|&}�����>��\��9_�U������ES�#_��/��螪��߬�_�c�������w���J��=��7��|�����J?��-��������DϠP����?[�~YO�w�g����-G�s��V�x�T���{�s���s���T��o���ғ������M���4�v���U���@�O�_����X��{?G�%>'����m~�b6m���f1�|B������Ǿl����|����'<���#����D�����<���}��w��Ṣ_����z��y̎=���_��/�~>~@����t.I��=�P����֣vD��>� �;��!;��A]��g���}[P�f{u�=��ݛ�ڮ��=�X���n��v��d����Ҏu�l��hzs�Vۮs^߰�v��ݪ{W4�Tڱ�{m�{e�F{u�&{q�Z{~�{q�:{c���㡇�����6�K6��{a�:{���ϯ�h��m�m�j/Q�um���e��Q��o�v�:�ݚ���-J�ۋ[���%�wz1xn�#�A�wzqzN/?�lx�^ȞݴYi��m��yX�l�?��s =�Au�Y��������:m�^����j��5��5*�i�=�r�=�z��a�*������<Q���V���%��wK�۳+�����K�6ڟV��gT�:�B��~�D��+Tn���to�;�zu��/�f����}�_��w�gG��]+|�kL8f��1V�o%��-v���|�u˖:��樓�;�(i������RG�-?Q�(�'�ZA��)�ҎX��/@%F�RG�P�+��������HI@*-)4���Yj���)m�k}ֆ��*k��*����
��-��!+)ȵ�^kkT��z��j��v)��fk|:����ͺ���i����鰱����s��V_���������lkLI���ǭ��!Kc�%������Ov�g��3�Z/Zܟ^�]?���}���g,NP���?��?����o���������������*���m�/~e�����0U:�_��S�	�/�~�[;�g��s�~���ԯ��/�������W���<m�����{^�k��tE�������*?hi��[=}ت�Jﷴ�;���vS��E��<�t�$����[���v��j�c�~���ÿ���s��_�ӵO�Yұ}jm�����l�/~io�䧶C�l����d��_؛J;�_�뿞��z�{U߮_<e;Tf����?������kھ��+�c{�?����C������+��ڿK��S=�tޛ���hz�?����?�����g�h-)�Q_�R�}��m��؟I��|<�M��>��N�ا��訽��c�ٞ_���^x�v������������������f�^w�>w���~�������W�{U�#����<������w�k���w�����Ǻ'�7��奔N�I�e���ۡ�-��lw��{��8���k���Kz�u���v��?Y�~��^y��w����K/�ї_�t�g��m
��m
��Uz9({b�vKܹSi�%��������Ǣ���i�o(��]m~Cm|����;Q��{�B��uI�o�iqJ�;v�	]+a�n�W�S����1�ï�l�_|��YĨ'v�V�e�vZ�:�uO	�ߴ#/?o�^|�b^z�?�[�{�K��{^�������);�ǧ�𳿴�����Y���_��ol����b^���xI���?��o������g~�sk���������W�1/>m�/ɦHQV]GT��gc	�>k��3;��}F��O��b����=e1��ڒ_�Ҷ?o�ڦ������e�|�r��fY�_��}�[ΞW-k�K��_@о�C;���.+8��*�ﳪ�V�p�꓎Xٱ�֜ceGwYE�n�O<(�z�ZҏZ��J�1�Dj'w��V��L�Z[f�5��\]�-/ɚ�23�J�X��%xْ��$��3���	LE	{�*C��ZN\��ʕ��J��Z�e��z������tB J��$k+O���lk.K�Κk�ʴ��B�mȏ|��%:ۛDa�%' yj�����)���:��˲�ǭ���z:ۭ��1��h���A�U�ͺ�n��G�޾NO}�]�?�mC=6�41:b�2,S'O�)m�������2�..��j)����p;0hgF�l������m���N�s��ԴoO�����J�Ƨ���S��Ymi�Օ��5%�J\3��J};>0doM���:��ؤ�5��&'=q���Azkj*H��ʏ�;ӧ��ӧ�ʽ}�}��{���oۧ|`�O>5#}���g�_����E,��g��?���}�������{�*�����w�����*��{�ۇ��o�e���}��>����w挽����{o)����w����{��!}����#����k���hz��9{��Y;��0>0��Ѡ���~���n����J����w�kS'mllXi��ǆlb|�������h��&�'lJiZ�̙S696j��C6����`51<lCC6�����M�7C�E�ߙ�956f��=���i�䄝���t��);w洝���<���L����sQ��-���ۿMo�;z;���y����?���X���.��?l�>�����?�'�|���/�>�o��l?�o�~�����n
��m�{eI���>M�+M��{�D�s����µ�N��=�}s�x&�~���)�������>��}���w�O?����}xn�ޟ��c���D����F;5�b�����`��j���z}����v;?���N��P����[C���x�Mt��HK�M��Z}�����ps��sReFZ��@�����wG���x��&:k�O�P~���N��i[d�m�N��h�z�MvU+��i���@�����������z����dk��w�
C���Wx��g��@m+���B;�Vl��%6ؔguqR1�,���V�~�r�r��RA%��v;��3V�c�y'�6��Udt�Y��W-��v��bU&��N�?b��&/�aS��x�}V�+ ���D������Q�������t��s(�����\ Х@B-��.���)����V�a�R|�1��(5�@!uH!uu6@��zI��Rߥ@R"߯7������R��@Eq��efXE���~�`�����Ĩ�3F��Ԥ�ilp0Zn�N# !��Ιs������%mɏ�Xui���T^u1U\LUS�zZ���o�YA���g�3�S[��tN�a����[چ鼠ıs���"�/���g����%�%��G&�ϟ�d�H��>��O>�>w0��O��O?�ӹ�"��V�,O�ë�'����P#�?uD�0���g�����:�u��=��S$����Ť�?�u��S@)P�#���;�~��)�`x�
B'�m�䐍���(0�	AiR0"ML,��*�O�z^�Ըo����Ȑ��ņ�O,���y8#�����ҹi}/J�;�r|_�u��{�-{��YO���{��+}���������J�@������@z���A4���R@�~����@.}����zn�0�P"��#�&>P9���K����������^z�Oȓ�ϔ�4}��?L��s����6q�%L�6�S�}���|8�:������y�_�?��뜾�v~\���fHF��m�����*lXۡ�
i���U�\f#2棝�6�U���:����l�����
�
d�ˬ�*��Dzjsm�[@о��|k+K�ޚ<�_!({]Uy�'B��\J@庪���&�FZKUV����8��F�.�5�\�m/wذR�l,�:�QWU���Z��廪���>O�,�1[0ʷ޺,+M�/5�z٪s�[^�.����ZʡW,a�F��S+����Y�R���/U�}�M��?��2��`gu�1V�mI2+����x�?�#������
���"M�ʱ��t�4�P\x$����߀D�0",���TZ\ೂ��r-��)U$0$@&�CRl{lPidd@Fh��z�����򳳬��LJ��Nɘ��[��SS6<4���q;szZ�JFN��|S}��TUؔ����!����o��[�;����7Zҩ�)���*/-յ�����%����^o*2Z�N�Q]g��I�No�g�����hz��9Oo�;+���U60`o٧M &7�7	zH��S��'�����_��M��_���K���>�H�ES����y�۶�X\H�<'O�}�{{����]�|���mX� ������.�1����0( 	VQ ��&��Hc�� ��q��Ԕ�4-E3��l\�[=�����4��o����y�w��u���V���>�{WpRz�])�(�<	*��O`��$ �s!J���|O羫-�}��w�2=��;����s��uh�I[�o�_A���p� �h����_
 P�ԏ�Cx�O��v�m�{��t�M�<���.�()��=�sg�bqvZP����!;}�ߦڥ���T�Do��T-8�ژ'���ʆe�OvT�dO�MtiXF~T��
!JJ�[ �ћ��hSq�UeS>[
F稞����pS��
*�Dj���nF�XGE�����B�VS �r���������2c�����Z[i����s���!)�����@����"�koZ~�n)�
����pP7��_���tA*]*)֚��XK;����
�;��v�k�Nu �Zm��JQIIUH��'t�H�%�\Y����d]#Á�^�e�����"WI� ���~�K�Ԭ�a���uı�?�
򳍙
����Q
��Q��%$u݇� ���f��,���\+��{:m��̨�ψޠO*MLMبތO�J%��c��������)��t�̴�����>�$h�
�tJoÍM�VRRb��V^Y���b���
R�Sm�ℌ�[~�iA��Y���9��Ӻ׋^3��"��p��`'���w$�6��O�>>�?4��
���P5s�9�B�8�)]
��k���K��ӱL!��[[�[ I���������sֿ���ax��R��P���M7:�H�ƴ\���X4�;�RD�<��N��)<6F9������oB�i~J��{q(��(��QFڢ���=�@:ooK)���۞�}_ �$���$���;������$һ2��&��M���B��-\�|h�/���ϗ�	ӥ��t)�>!�_�?��"���F!]�RxN4]Z��&�����.�#L���K�;�� F��� }_�%���)��K����:l��Ŧ�l���PFRLcR>@	U4�Z�J	��
X�R(�ͥ���J����l��d[����VIU�
H�:����d�HU \u���J�/���pY���A� Ȅ@��<|B�/엢]�	���Pu�Kq ή�L� �mI��=��J�8��j{y��$Q�z�2�ow�Zki�C��<՚-7v�U�lE�!K=𒕥t �*���:�8�j,J�r	�fU����[=`�V���ΪWo��)�A�>AT)�n���ҥ@����:
���!`���ؗ�`�p�+��"�0rH�w�R��������ɰƖF�#c2(�ԣ��a�Q�G�ǵOFkj�&eH�yS־�.�йmRd����d|Hӂ����:&I���[)�m��v��Zai��WWYiE��U�~1�?LJ}����;%�M+���:}^u�?�t:z����32~jo���n!C��7pW�gRI�J��G ���;���.�ӡK@s)d�o�h�N�h�@ɯ���M��]� Q��ϟ|doKQ ��z��
|F� ��$ �q}�$@*�I��mr��:�ɡ��wM�o��߃�&�$�ˊ�}Wo	@�D�ο}N鼽��x[0���0�#��ݏ޳����҇JR02���w�T4]�/����B
t)h�{�H_���@����3)��M���K�߭�H���M��~��g=돕>�z}��z���(�~�Q��ls�4u��O
iL�(���*I�1�(���r����8f�z�?�[����R�R)������ɐ@C��"C@ʓ��vX��
B�R��U�H�J�R�S�@W۸.�H�� 	�P���5�
�c}��:G��5��r�Ϸ�Ľ���՝H����.K?t��'T3uNn̛V&`���Ľ�(: �PHm%z��3���:�D�7.� DA� ����L.��}P�/0E� �DH��'>K1Ej"�υľ0�eHmM����Hc}u$+35��|"R]]��j��F���PD����WG2�R#ٹ������pd��Pdpd0"E�F�=��D���Yid��I�'=���),-�����G�ę)O�g�#���DN�?�Ϟ?w62>=�sK"N$;?/RRU)���J�*/����HckK����#��OE����F�T�ԹS����kN��~%Ɉ�9}z:"��"z#��?{:��[�#�A��?��_>����B�q��>�$y��	�g��S��D>Q=��������ȧچI*+"�xd<���\Ү�?������'��9"E����ȹw�G�V"R�)2<<��`䤒�QD`R�F���"��'�����hD �4>9�<IE��|;F>�ƧT����߃���7�}7|O����v:�Μ'���{�\�l4���8��[A���;r>���������������U�.���ςх$�xd�n
��>����kyd�/$��B��[|.$��I��ti]���qi����k{�>��}�(�>�P��w#��V��"��LD�M�E���n�L��G�["}���*O��������H{yd��62�]n+Ӿ����U�Q����G���#c:�^������F�{j"�~�0"���V�*�W��ꭌtT�E��?#�Z��Ɍ��f����"���Ps��$ i[�"RK)�H_C~䤮;�Y�c�)��@�ڊ+/�~���]��\';2А�ˊ����c��/Ejrc"R�:'F�#��qA$�~�u�mK�F�ڼ�H�ʕ��d��H?I��BD��4�G�HsaB��$9R�~$�X�i/ψ���E���#ME�ڗ��N��R����4�%ןg{EF�_��k��ꞇ��"�_s>�^ +��    IEND�B`�PK   2acX�#�(~ I� /   images/e51fe3aa-205e-4659-a3a1-ad304791dd1d.png仅W�Q��=�!�C��tI)��t�4���H���J�t�tIJ��Cw���>�z�ᛵ\�f�k���y����	S�$��N�����TA _�*2�X�����(������BqO7x��UZ�U�����������拽������g��#2�$/�^�q���~�(~<�}�̨_�286
�=�<jD@ �G��a�nm���&lz��p~�r�а,��b�I��MY!N�HGO�k�/Ɯ���c�ܪ����E����)��U<�cO�v��η<zyt$ǞUr��zĽ
�!���D���h�r�0��jc������`Bw��d{���V~i�;<�٬R]E�Y���z���kWA��}l���3���gӏ�x����\����	�$	m�u)�Hy����@o>����t"�o'�������^1k�!��g�l�BH"\b߽�~�����1��O4х�bs���_�ч̜�Xc�2���kN#�Q=��
�#�[�e�Gl��V���"�#�Ü����fɬόzP3��hyz)�*YAPW/��	�V]I����')G6��������\ys+)��������R��F�|>�kb����p��pdG�E3���g�}���|k>{C�����8a��-.����06�<�t�y[謤���<I��#8	1L��C�~���@
�Fʩm3�9�oa�Vi��2F+J���K]����ԟ�K�a]je��Պ��}+O?M�C�P/Z/��o�fs'gDDmE��h&�1�^ۗv<��Ԟ��)�F��3�}���A�gP��w��`�y�]5;;/�)��l�(֌KKϩ�I� ����c^�{��&���ar�;:��nż5�#��ݠ�������a��3�v�0�s�� �\�'��Z��&�_EE@ַ��j+^/���_E�9��R����]�O=Rf�u�2­5��r�J����-y�&e��=��&��c`�G/��QZӌ��Ablz�k�7gU_2����@G�\�ل���߁�@�o�^N�y5w]�����l�~�M���X�:s�O*��qǁ�/m�3:P�X;�xI 2��r7���*i
~�W˲����͹�N5����<�Փ/W{U�����>�kv�$��IwU�.�)��M��6�c{���mR���H�����c���ʒl���&�}��<*ޑB;��ϑ���>g�.T�|�"���%��H�
ӦD�� zY���}���a���H<QZ@Ũȴ�w!/���?s)j�͒oa]x��oFh,������1af|~��K&�Dz�=Jߜ/N�m�ס�c��R�+��g/e�|�Vhck���y�f_�� �X�Z��酳	�����a���z��0;%0��ԡ�mXbp��r�8�?��u8�gvܑ0	��6����a��ԻGO%s��0��sv� .��@s��Z��=����;R�?� �=I�v�V�0|�褣��I��k��Q�nm)>sV�N��u��r5��Z�J�����Mk�p��I%#��F\�o�(��4P�1FO�3����׊T�@w4�9�VW�U?8lX���3�ί��-m�C��Zb�Ԯ1�k�0w�_m ��nq�%����$F�LO��m1�"�~4����:M��_N�׌v�>��_�	��7�z��N3-���Ъ �mAHɏ%uhw�	����LF[�,:;���	�����chbe;%Y��J$���0����G���Zi�Ȟ�m��_��N��3�V�1��xN_�ʋ��:p���=���`�&�3f�8ۢaN�U��e�s����;�8h��&~P���W��_%v��,��%S��b��X��࣯��]����������u�
�P>R�Bp��)�]�	���O���tQ����>�W948����b��R�<tL+�88�WFJv=��A؇ռ����]9ޘ�%H��P��	:}�0�~�n��5])}�%0Nļ�e�qC���.i���M�[�xqq��\}'f����V�wd�O_g�^�"/�>��� ���Z�flȿ��(�d�e��k�7��캆PR,9���\F�x(
˟�����8'��}�y��%��e�W����l�H("
,��'�MJ~[_�����"�"���Г?\�.�5H;J'BP�e�
}G�
ՠ�D�˽���%bآ�"�d�����8?�p������'����p������G�󇻰�0��9��1R�����`)������ �2[�J�6��k�~�g��իD��#���I��S��oHm���In�[!>��[1�p_;��>XBC�x���if��nrԺ*n.&$��F2H����،���a�Ǆ:j���?H��裡�e�w��X'�U��@vN�	vG�,s*eR��c��R����f���]R��C��X
<86M�1�'�=v}dz�b����Z<~�Ƶ��Jz#���+r�c�><�$�$f�w/���B�O����iԚj}2�.6��z��I���X�$^��W4�z�yb�~1�C�Nu|q�2��bBh�v�>��h�a�M�Ʊ_W#��fc���)�������'9��q��v�8L�d7�7:ƕ�d�S޴���Jw��\�����X�����7K�H�0T�����ታ���`<���H����蕓F��4)=�/�_�}g������f;���f��>)�:�Ü����Uv���<|�/��Y�L}+��ԛ�ѦV��Xϸ�8D�SZMO���(/W�[��췅W�F=�;�
`=�]k^aw�&���|�Pƕ)������L�Y�Ğ�xj���<��_�*���$���"B��b�Q�W��	���>�u�3��	�ث�P0!������K�4��[�L.a~|C�Q㙞�2��[�w��T�wCV����EMW?^%��<��5�sU���ߩx��Ʀ��H(�O����R�;k'�_&�>y�݄�Z�{~`��"4@����Mz��ۿ>���1=X��n�����I���*!��]6�u$t�1�oM�${���w����cR��{��#p._�ɋΓ���k�ӱq�E��=[s.�� \ܕ]�I��8������<�iz�������ճ��)<Z�:�Eu@��6��51���K|;�2v9|�x9������>h�l�Aԗ�?����y�t,t���tN5�Nk9�l����+�����0�'��p��$V�u�Rm)}�؂�0C���b�;Tz9��5�EQ�6�+�y�~�����V�"����o�q��5��|��"���>w�j݉PZ��S�FP�??��Y��T����aJ����:#�Θ=˓(��-v4����Y�oBWQ\�"?��5������7O��PP���t�,�ݏJ(�Wẁ������n}xɹ�g�_��=2�����E`˃����H��n�!4g~n�����Sɍ3�%d�"��EpӒ��:��Q���Q\1=��h��+���nM`V��g^h�4�i�&z}���)epzl�7mS�<���^�vG*-�t"�.k܇0������ٮWW��B@�����|��B~�-s�*�<o���E���f�^���xi��F��s��M ���òB�߯��4�}p5�=H蒑�J
Æ�ѼB�^���{1�%���8Ʉd�&�K^��g��1X{���p:q�b�(����<��N,���Q�t�ڔ;��I�'0cbMG�Y�¢�Y��C�U�%��BKȴ8�6�W�� S�$���{�/M?�1��˴U�v�׍��O��������߆�&P�6<�M���և�g�Ϻ� G6��%$yᘤ�C�;�^(��N��Wv�vZr���'�GāHH��L3�[�VT�W��D@2�	�h�˓�pΌ�6~�����XB������@�k�="��v��;��h�\4�:��ƫ��U����X4�0}��C}x��G�����9Ǿ���O-$��xɑ��H�?L�z�� A,�[;]S�N5|윱��);���@��ھ�6UG���X���
��fb����6l���߫AB�C��H�QZ��l�Ccε荹bؤ�K���e�8�2����9�O)��5��Q��|4+ytE"�O�:3�1ٚ��5�HۊyI��к��h�h&�̀'5�x ��1�f֘ܖ�Ia�~��f��7t��V��q��|�eU����k�،��*�[�}���ݛds���5Gn�q��t�.c�h��W�.�,v�Za/�"hv(��໐�2���be�"Q�l���V_x�=��Gv]Η?�@��28(l4�����j�>Ki�f���.�Z��C0opbcҾF�5�v����z尷>˪��a�Æ���<�W���3e	�ֈ�����{G��ct�b��ٔ����kQ6����pĝ��ia��T5���|���n:�}z~�wz����6�
`��>bqi 6Z%�X�V�<cOQ��/�NkϜ�ZZ�Aaic��&��1c���2�b�y٫���pX?��p�%%�/�E�z�D�]?�\��Q2�?Lg-W������-Y�۸U���E���Fu2
2Bd���:bͅ����eDVL�F��˸?��؃�r�e�lU��u��|o���q�̄ǹV�1O�������qB(��cT@ݮ��slhB�N� j�x4�쐈~��ZݷN;6���P�P
N���6�6���ػ��MY!��f�Y9GH��+E2,��ў���''�����~Yt�x0��w}�WN<�-�"$b��o��ҍ�j��&��V�|N��i:e5IM���J�����Oo��e��F� �p�׼(S[S+<ɗw��(���Ý%�~sn�K����ڔ�d�'ϽG0ñ�U�a�����+n�u����K�;:�b#4��MG^��`�?�����isӬц���w���]{�vz7��h���ټ%s�o�����٨8����GdE����c߻�=�N��.�>~b�UD�)�؎�.z�)ܛR�s��[���BX����m�["�G�h�=ҭh�s�o$��~�Q�B�٢�
'YLi{�@`W��	t-qk=��m�JR�٣�jB���/JQ�B���!����<�������55�k��O��͇�圣17^��|g��U-ote��Q��y����z'6�;�$k�L�"�ʘ�(���VJ��M2�6��)�;<kE)��p����cz�DaW� 3ǡ���,��#VH�5"E������H_���ޚQ�_A1����ǌ��4u��2yE���"�kM�V���N�ECn����@|�{}��Mo��B��LcN��P��Xp�W�7W��O{���/�4��U�nQZz��׈>����'
�w7�� ��|F �i�����o��s��q,�� �)e��p�]���y�5�犬�����u��֮X)������U>"d�$��Q8��T+� Yn]Z�u�c����er,���MZ @�9��~�d~����V��l5H�̲Ng�����U���a��y��cK9c
w/�B&(U�~،����	_����:�\F�6yUJlC�;>��w�����!K:E�D�(T���=C�k��T,U����Z�l�V�Ƅ)�5�԰�T�T5�M/?a� �z܆��Wx�~1���K�]f�H�nElO�5,���I9b��iu�5?t,q����r�{�؈��{fR0�ԑ��/��A�`��5�_�Uv�@��rP�I��}��N X���e�GVJ�p�#��fO~_�1ܟv�������������r
��Z�p�7;��������s�!nl�l�6�;.���04��'Ⱥ�^G'��qd����*]>�ډ�%f��6;攑��Ǐ��K���L� r�o�q�K4
��3I��#��I*k�2��$t���R�u�H_F=�H���f�heq�?����>K����;fzX�T&\���w��P���۴�eWg�ŃM�l,�_eSӿ�kZ�PGą̃A���z�;������S�P]<'+��7�5�ɲӧ%��PHf�0D�������l(�Ga_���v4�ZtN�hio)0����?������mfޞ�����"Y��o��7''�<J�X1޵�����AXE��?��鉷*��b��3Y}jw�Z_��2e;اК�^!^�"���A���W��a;�R΃�5¿�n�(��?���J�g�S�ו�`]�t�]6�B�/JNk�V���d����C?���*o"űZ�v`�.��f�%�=���u��S��r�6�T���� Gs��LNW�ig˞e��3�&��.�YWﭭ�r_�	�H�(�a_�eC�xPtJ�x뷭]	�rX����������1�Ct:?Fqdw:��\�d����*i'_x�\�"��6�-CJ�m�}��
䫃f2=��5���F���p�����n�Ѥ�J�\Kl���H>�|�ֺn��;�b?��!��c�3�C��h.Pc�c��Z'�Z�1�v� ̽�'�!h��C�����F�BVC'�=��y��f���b�b�) ����QB^j�eߝ]�>��{�?:�&ty��]u�EĞ!`6�"|�̑'��p*=�w0���k�+a3��E�d�T���z�U�|_��nU��\	ED�)�a��g����� �L�8'h?R�����e���0���`bz��s�|��Q���tx�=��EP'���x�ph�@��e[����4q���LN��!�
�z�6&�6Ǘ��t�mp�;nB����[�1�5s�R�5�-7�sl�P.�'n�m�rXl���7���=,/�
;�2`fW+Bn��u�m�RWB�;/G�H��5_Q2�i�[bD��bc(��B>������e2G{B~w�fOK��3\=ő��L8���xK�B�D?�&fwy�d�_�Ue�Hh�W�+N>�e��yZ�E d�d�<r��^ݠ�8��Y��u`�i���#l�P��mB�xp7We�L���@M�6�kUf���Z[MH�tA(�g���K�EG���=<�e�.N�!�nϙ!����L����I�X���c��uO3�)p��.�1$�ɰjc�T���B����+*4����q�Z�Z��m+Kr-�L�v7q����������Q��_o�����Ǐ1��u7]�uz��:���_*���+�A�c���s��F-���N� e�T�8����`�Ub��^�v�f�x���l�V>���t^�ݡ*5�Xd�m���g�ci|p��g��ⵡ�PG-Q�Γ�Bs"5���M$))�0zyw�;Ɨ}&���T����u�2{ŏ��(9��z�ޖ�eɚ�a��Ҫ�4L��QV�X#E��v�du�� p��r�⽠oT[8�z=%l%"{t}�2���+�j?-����w�޳��=_�{`�h¥�^hU����,����T��F
:����M��5���/��n:Ɨ/A����C�&�Y�p�(���b�R�o[�b�źwQP9�1�v�X������ә��`�E�������-����^#��I�#���N.�������R�w�`]�̅��ѓwDh"��-H+�
��s1��7mA.o��d'���𽌨UR�c<}~�kC�y��5��L����bh��߷�&ԅl/�DYtK�$JDg�ʦG��g��H�qH���8;.�T�\�3}.�H��������Y2_�LV�+���a	��ä0�Rf�0�+d����Ko�m}ױ��np�����DR+�v�j3�����Y����q�h��w+d��j��ҩ8�?#���p��+�c$��xѿ�<��6�Тڌ���6joy��֠���Z��z�x!�>I)^��HJ @|];�ͤ��[��[y�_{^�t,Oj��z(�W���J\�Pns��n�������4ZlV�Le�X�Q����a�Ox�KUy�p!�
��s&�����z�UM�&�jz�Z|�b�?�]���ι`���ú ;�a�g��]�#_�s]���yE�m(��2���.����[�/~�j�#a0���o��XO�Ix��.���v��[����?���0��Zí���g7��5�l(T��l�z��T���s�Ee�p|�Y�zxF�7#?��_[���bD��=�ѽvȍ/K��絡è���Hx���h�E�����t_�rk��R�9֡�I?1(�odo�^�^#:��ї��lC�Z�*��,U��}̾�C���Ս�6qsl��-��!�ۏ���t��$Y��9E��_�4�%<,]�#F�F����d�}����x(�?:S�݈Иʪ��
Q(�_(�,/����De���^�ԑ�-%Ev�0�P��ļ����a͈5͟��tG�b�hql�fb����������d�.��^�~Y��-��E��5a��ɝ�7*+v6��9k�����i�̦R��W����8��&j}�*��$;,Z�%IO����A5�W��b-15C3��(@$Pt��eĒ=Gō" ZI���YV�SB��=k�2@�]��Fǿ����ɍ14�;4������L���j��<b���|Yc�$�N�.K/m�EmBZ@�`'�p����>sc>������j=`[���D����d��~��Tt5������L���"��X�"p#�WV$q�}̆z��<��	�RB�n�U����'�q���X���;r�if d�ډ���P����#����%썺���TJW8���+�t�ڋA��L�!=��S�K9�5���4�E�M�O�J�y(�#�j���}#!h���������{,t͇�x؟�E�,�~�'z�C�W�:v��Դ�N2�F���э���<�ޙ���� i�S��-*�4z-�n������RW��2J�J���Ɯk@��N/�Qӏ=�l{ ��=�!�S*�-�Q�p�J�-����B�晏��q���ow/�k��P�t]ᅂ�;@qRl��s	�������⢝�%fcE�g_���;3�/.?���x��;>��k`��{������ϛ�M,_�@��c�����o��g�֬�*���6W��&+酔v�L�U��q�Q5�c٪�Yh�Ľ��+���0kV�˃�%V��ѷ�'���^�ھ���'�z)����#��b��ױ��`g!fتj�ŷ�Wvr#}$K~��U��MeN�,~S7�S�'���Gs�y�����:�/�To����$�m[�Æd�������J~��� _{f�#,�p*��$z�D6���-.��JϿȹ�+����BU�D���7�_r�3K�!�ͪۍ>����w��e2'^�۷�-�Uʅw�*�+'���葼���`B?D��Z�{i���y^(�cw/�^�Ghd�K��V�
�C;�Y�ʺ^���y��y~,�PH���e��OP�U=m�q�]��-�!�h#��+������X� �����'�=���I�F���"�k��Xt4d����5�'%m_�W�%f�ϙu�*���|�t|�]�{��o�t򏙉��Z���qk��dGri��k��͂o��ihg�h\3Ʈn6��S��q 	Z2!��¥-˼c{4��,������~�)�j?�j��eE�����C%�����z��X��K���mb���/Ճ��i������c�}v��݋�C������U�VD�"����?�~�3 �wɉ)��p�c�>��-���txl�E='[:$��bs#���J�;3LM�	��J��F�3)9�3H1Hh�H�M�!#rg�"�BX+��,���
��T�M��K&�QzY�E����|nhL�A1����#�@��*�3�"���9�����|EL��ҫ���	���G�8��l�^N;��R_�911I�Æ�kר�.���D����8�Q��㾁[�s�[e�jȯ�p9�>�-S�y��zű�-�7�}���b^۵�m������/̊C�a��*��n�U�R�<Q�gDK�A��E�� �Խ$\[��sjY�q���z(�:�;��	-�L���R�N-=-��	����(��!P�|�������s�\�W6*n�x��a�#q%�$}�2^:|�z��Q`釋�oaRZa��$݃�!w�c��[�����4Ծ��{GXB��],;P�;-������k�Ʀ���]lB�Q;C����ov�x��=���:�E�p�}����N[����˾��{{��Lfˇ�o��F��dzdۿ?֠��l������/H+Z	���iYa��:3�@'Gw΃��C"�B� H* ���t�OR�0Z�m�R����^t�
a[�!�؍j���ڻ%�D��Gl _��^'r�����c�_6�W8�_;��Xk�S� �K}�V�qg!,��=+�"}*���c���C89���eduz�_��z��E���CC֤��b/����y��9>=R�r�9�ܪ%�.�����=���o}�����
�d>2�L'z����� �'�������ǁ鹞��踜�&���b�T�plb�NĴ:�ё�K�<+a�(EUGf!z������r�Y����:2z��.�7 �B/K�:�]�5DkiסL����b��K���s������h����o
��e"J�O�:Ѱ����`-������T�I�s/�՘ypx�9�:�%`Nz����kN��G�qz�P�9af~�#gpؚ	��G$���(�O�vH��d#���T��CW ������5������(SkHP�dN�U��Z8����;�l�?���@����ª.��G��J�)�����m��߂�|9�]�f�*&�]r�JĴ�Ҷ�@��xPM����3��#o������9���$%d~�� k�DB]Jʾ�ۖw��au��۬f�qօ]��ߢr<�,@d�ʪ��ڔ,J�ʟ����{f냵�|��FH�?�D��y��ĆP*Y�9gZA�T��ׁ��r��B|��	�%|�8��iЋ�f�i��c�P:��.��;lP�Fi�TF�w����������đ�1Z�{��o�4�,L�-�\)���[�,I @A
̘�ޕ�R��'�_d�����[_�g$�plWc�rd�)���Ƒ3h;����]�5]��������.m��&�U�n�m'�Ǚ�f���u�/����q%B�DS��T�#�}A�&g��Q�Wj�އ������j�j�����&}�'BS�7�E� (��J��yfgӯ�Ih���k���z�Ui�-��mڢ��tj�퐟D��\�S����,���q�,0��؜�<,ͪ7��>O�I.�#�ɮ1��ٝ���8k��A`��i ��<��5���v���>��|��/P�/�w0l=j�}�#�*?<��+C�h����3'�C��%�G4y�X�bW��U�0���AM7�qņ�c�9�o���q����"��׽F7������ݳ�W/��(J�#� v����)�S7ir��u�$,��k��4�G�·�f�����P��z᱉I��Z;Q0d��EVJj���-��^������ �f�������˹��ª?pS��>[+c_	�/�)_�%�>�#��������n���s��*P��R�����އ��ќ�#�� ����l����8�����1ȥXE��8���$��F�����L�ws0�,��o���yl=o7y|9��+��c��X�Y�~�u"����A�e����T��EJ�M!y��hݽb�1��Ϯ�b�TRGaZ�W�%�t�����gx9ls�7flڳ�k��y��ŝf�̪�C���6�0E���Q�Z�$3���	��a��k���;�]{�MG�A��ݒ	�1a��He����=z"J*-�X�6�{^���P�Ui\�5!�uz���Q�s���ν�)�h�{��i�U<��}g��^|>eY�?0-( H�y��ظQ֚�A�����-��+Ƴ-a}���qmR�� {�=0
V��_�m��{貙��v�h�ngGM�Db�a�_K@�4����u/�6���_����U�A�$�As�j��T�<H��q�$�4� r�0׺����z�K����o+�(a&�L#��Q(,����@`G�� �/tQ{{����PH���J����9Wy
��' �` �Is�M�{���~�e�X\�9�j�6G��iWHޠ�� J�S{�⊗*N�Y�����H�N���OT0�j0q�?�d�h��H�;g�N!�}���5S�G�Z��c�e�`AM��l�?iE&���Xʜ��<��X��\�s3 lJ�3���ޕ|��S���ta�J���5s��_��g���l�5Y��U?ݱXg�L�p
`v]���d�5�?�=#*�"��n��KVÒ)��,���-�E�6�Q����|v�<:0�y�誉m��uݑ��G5��s� �r��L;��5����
�J���IAm��t�L��Qe�p�P��g����Ţ�B+$��Й��O��Z=dlK � `��J]��OrԵ
��%?^����+�'��6`����xD@j�N������6`<�,�)���
~�H?o���,M���@�(8aF7��QSk��z�^z���gJי�O�ي���5�c�I-�b�_�k���m)��&�o27���x�$�^X{�tjR�:�������T���-�����d�� ���3���P���M�f�As2N�"��hV���_��pn��+�Jo/Z������$/!��#(�zi�#�$��8�G,�AC�*ӈ#�}2���Ĉ�5��a}�zL>��H]<�.F:�:�Y�֑�ѷ�Pk������&ͻw�s�TZN��p�����-�uW�	UC�j^�Ⱥh�M�遴��ȒQ���G��;�����7���$U�_�K�&�y����dqj9J�gsHy#��Dkox?_�]�Gc
�d����aWZZ��9�X*X͖禸� ��~c���{P^��KV�P��Jǋ��}��9�ɴ����a�x68G���3Y�#�D�[����l��a~wg�3.̈́��qz��cg�+�Qk�������3%�B��a��� ��EW����6c� ��r�Z����y�y�1->=`�ӵ_&�s12�=�%�_1A�#?�)���p�m�L�B@pp3�p��E�Ka�b�D��̕�0�$��c�K���\�.t1�E�����m�"v}�`�<���z��zQ4r�B�����I�5){�֫q����^	�,l(��&��*Z��������:��ԗ�sz�Fr�,�6�~�\[����%�I����������4+�˵�t�$�>ZВ] ���7����e�5����{h���M��:����Io�WvC��_��i��1�%&`��O=g�Rȡ.k!�{��E�!�?j�c�J�LVF��j�|~��\����39
c�oեXˍ��f]�BDoI�W�������
�,���N�8<<8?{��iA!`�W=�_�pT��.����眛���82�p��vI.�v�HB�8��<ZoϹuz[��r4Ű�P�5��|j]�&<���z3~��X�}9�[寵it���32�!3����DB5�B��D���j��
��HT�߶l��Ю&a�x���AQ,|��A���$�!W���!0��b��肷pe�H�*�u�M�h��wLҟ�Ą�߃��i8�^�>�O����Y3��^�Հ��G;u,%����6��>j4d�E�c��+ȇSӯ�������A����1Ţ�=!�MK��<e�ﶆ� $UK4(�v�K�O�25|
��z��Z�ԩw�ۤ�痃������)V�E���a
��䌷���u=gF������v����6ka�E/�BXW�s.)O�K�������k�?��g~��t�=�{�qw��L_���&R�S����W�u�΄ef0�Ժ��p�ހ�C�S������ �t�38[s��\��{/��^��+����L�7��f���X�|HΌ�>S��?�Ŭy�'�%���U򷞢l�Z�.�ǽ�/.�$��~�7�a�k��@V;�r�hW���S�d�n��nn
	�Ġ�x��I����<�f��� �W��C�
RR#�ۭ"�����O2�GY�s�
�_�*w����/L��Z��&ɘ��=�N�3Rm1L6��W����96�� Bƭ񾲀=���m�Ka;6�Ź˛�fa�H޶�~a��-r���54>�����F3�Y�O�@���g����Q]cۇ٭ۦ&u�H.᷒�WǟFT��?���{�7Πp�o��_s�m�.7x&5P�n#����q#�&�Z�|�R�C'����7�.�則��?�F�TZ��g_(o���)t�/����0�wx��P�[˘���[�J���GM�����w׸��ȳ��o��J6�]�v7Ǐ�S����h�lE��Іs��S�^��_ޙ!9�0?���*^���V��PG�/�;*����a0[~zP�~����?_�S�؟Ɯ�6��a�ڛvb�IU���[�m#h�(�D��;b���#0�4�GB�\�[d���aݺ�lA��ō��oE�K>l�~7_~��f
��e��������G�u8!��ٍڴ1���ă���3GŻ��I�����M#Zڂx��e�'�d��k� ��ue�l������Y^�N �C6����H��G.[�1@sT`����2����D��K�������ĠX�b����&�|�~4$��r�ia訓?{\��l��),�"�Ȇ1�CO��2y�l�O�L�\02�I�װ����+��@4ޞ9��A�i���{bc.|�%�7J��f16]�� f�ʀ�?&�]˵��I��$ϓ��g E=WI~�$�&��aXs(�J\��x���F!�~��C�zkv	��������O�oSmR��<Tl�IG�ݲ��_!�Z"��9%/��o�4y�⩴�_�	'Cy�ק����c��wmlE �0|f4"�'�;�%��������űl��Y:U�}�sfX;垲�y��qq�FACJ�_3�l��~(���?:�@�4�4��T1�+6rc����po�jJTQ� ���n�K,7v���[���=zl-�Ə?�0K�j�H��>���n����}93:&L�G�������brj޵��>�M�^���:N:/<��ǖ�#�~�gX
�&	�5�*qti���GY�%~��+���g�p������9���Nn�}�ޗ�/�2��rg6Oq�_C ̺��</�G�%��-�{�'�XraR�J�W��D��b��k]��E-
HQ��f�8p��Uz�'wt����o��a��0E,Ȭ�� ?��s���ւc~	xp$ֲ�쵘2����Vz�U4�1�[����	U�O�����T^~4 ��r���f�J��~@Zنf]TZ����x�&.�8(ǅ����pʚ[�
��F�]DK����7jv/;-ظ�������#h�U�R�? d$�x�$�����>�G��j�}��Fе-�$��;̝��	+�'&�[��H 6(�i��{a(����.�W�D�����i[�}�n����wn��2m�k+�2ٍ���^:v��'���k�C���3�x@Rc�}Ҟ��Z;�L��G3��J��Oh���y���f�8ƾ���:|���/+��[pG�[�Of��?C�ǧ�pţu�w�����,�&�����_X	˔0�{�=m��e�C־p��[�C��C��ow�;XpH�7����LZ��MZ���F9���R1S�n5=x?km�}�&PTD�:l���No8���"|�
��żn��ĺ�������P�f�����By?r����v��B�GhY�lio�(J�(�Kzߦ�8�"m#`�WM$��:>uKs~\F�_P�W۵�	'�[�3�0����ň�v,�iǇ��A��c>O���,L�ҏF��Q%u�_�m1�o�Qb��W���i�ITq�-Ù�4�(P���Fo�~aX�4����!���$l����"O|��E�ɲ���7z�Q'"`��O)M�􄩊��E�Ps�Q��k��4 �f�=_�G�Y?�2?
i��6<�A����%$��qaT�r�����_������Y�3%@2@�sCԯ���.u�֢�^�|@I�Gv���~�ms��qz�5- $�(�ן#� jfA"�%B�ٟZ�G��'��k%�Z&�fM�|������%pn+.�f�>�斑1!��؆-�T�ܶ<2*���֭�׏F;�v�(��-5��x� ����\��S9���W�ݯo��;4�T�d�11AMz�YJ���S7�v��}�%��?�fa�I�Fݚ�]��E#���\���ȡl���p����ǚc?����~��/X��R61��'�h1��Z�~T}�.պ>��O�f�|2d�x�[ҍ1���fO�`�6�c�/���'��RR/̾d)VZu!�j��� �h�V��X��R�ʍr���8L���(Եr��=����~+��f�S�fɬˮA�oiaRE�8~�K%�9���l�VpjT�12�w/b��ed�S�E����p{�2�?�{�|Yğ^���`.�ׁ�V%f��;r����GH9,xyLYiN�M[5��%��_[�Q��E�a�~rEv6�koi(��\��쇝os���.&yE�Mg��3���8��.T�ơ���]�:�%י�)!
kz� w ���Ҟ�J$atu����E��W�����S�jK�.M��������������Q$8www.��ww'�C�;!�Ӹ�C���ws�}�8��h�w�%s�Y{U��E���[ϴ�	�E4��z ����!�|ݰw��]��)��Z�;Fm���gk:(+L���"�g�	��h8zQ�Ы���(d�����B �#&���wf&���ؿ�3T�X>,���U�7��Wf�y���g[�r^����"�8�2��7��)�d����3.IAx��������q�f��[��z��! ��+?�Z�e~l��\^9��~&�#ؘ"�M�R޳P�eM�^��H��_��8�G�t)�?�~02�p����������\˸Z�Q]~
A"�wyl���ڀ�w���W!����J�
��O��[���[.��A�%�� ���-�.�KV1�>��*�q��&��}�T�}`�^r�b��jચ�E��)(˵ �S����t�c����mM#�Ob���������pXa���>��G�|�+���@���<�g�k=���Z)�ۿ�N
��`��
㥙j��
����'IXENL<U�v��w���=#���)�D*��	�"e7{?;�ߪY�kN�FW���[��e�F%�F�r.��Zl1s�m�r�P�e�I��d2��2�P]�w�?�GF.FK��9L�?wZy|{<duo۲8�@�qY���oL�F\4���#q��D�[���S���su�?2��\���IKfl��~���gO-Ǹ��{��Y��r7�h�|po�|]|�U��FZMg�7����S�(sJ���IF�x�_�ixn����@˘��Z�|_��߈��B�s�[�ZP�4K�3�s�I����}��'���
����|�WBO�N1I����}�"�]�
}�^�L��o
u�҉W��.w2o��|�X"���<���?P@eս|Tf��o��?_��͕�ğd�A#��b�9Ѹ)e���J5gZu���V�aqp� A븈��=�ĳ��3�S�{+9Z\k���e~�������w{���� p_hޏ���3a� �M;�Ѐҁ8���R����p��|jŘ���զͻ����gau!�=����~�q�>�ى_����f/ʹ�U�ߴT��yba.��e��������dc���G�P����G�?jAg\x����,��,
W~�c��C��P��^����D�U�m�����_�/��:y�_�Qەw3"�n*�������Bv;�-
��(б��9̠��L��? {�0}v>�֡�xw��sȟ����m�ODO�dL�vkQ�lhk��b\Y��=��}]�~�o�9�I�1P�| �3�*��;���4�/��h��k6���o|Er��q�4����i�.����ۨ͏-����sI���D5�:U	���G͏�I\2�Er�`ե���<�f^�o}�oBmK|�e76=�&w�	={]C7|� ��̲����+9ҧ��(���q��V���@��;[:���E�4�i�A�K_0X��O>��3�QxvjZ��k��F�=�w��(�����y'8=	f�6���!���J�|�����g���'����q��K�k0"l0:Â/�����ʤ.��ֹO�,F)r��{�ւTs���K>���cUf�,�Z~9��r��j@�q@�%�K�I<�'= ��=�΂R����d��{~ �z����x+$l֑Ч�;����[�	mP�z�|#�&G�8k��������U�/�y����w�60���S��L�%�:����l��7ю-+�z�	2u�����}ib�Ы��[��k��k�$᳼��^
�{N+�hM�"�PQ|г��d�h�(^z乢^�������t��m<�f^�Ug�i9 �=�$��p��:'�h���'D��>W#V�ì��:�!��h��i� ǈ(�k���
K+|ki���ꆴ�[�dɵ����`�<��������E%�}��፳|�mS�LP(;��r�G��5�����ԁ]d�	+����ЖȰl��ul���Y\���N��P��383�n���B��>)s)C�fj����ص�������]v���h��S�iW�A�7���]�V�a��qooPZǬJߡ���1�@�/t��o		��ӏZ��x��g�L{����'�I�'͡���LO��&��(5�%����'�4�f�*��)a�	r��,�D��O�0% �|\�)+\��>������.IwhZ�y�5�61B����?5Ɏ�,���w�K]�������.�]��"W�N����~������)X_pܹ��a�]��R�Y����vý����e�Tˆ�q�EˬÏ�	6�K�5�?�5���{�l)?	5�����4��b�e��S�
{e�z�Ri��c����������r����k,���VM�����Zv1���*��U�V�π�z�k{���K����ӍX��֤+$�Ԍ�H�/�Ͷ{���S��F:�~c��A���F����Zt[O�)���tN��Xa��zO��͖�Aaz�R�W����GG8��x�U\J^��s���NR�}�3�'�8����Q��t�W��/�[�|b�.�j���}��!� (Z<˶q���� ^'צ���i��A�$���4��-Û�I��|�.VBS{ԫ̴��;V�} �\�(NX������^�2�RR5x)�� ��J��ﯪv˥d�v��?Y|�y�n���~�#����
)�x=%E�5J7���E3�_6Vmus!�]�_c�}Xz��^Ds��!kF��8�� d�U6��������G<=�WD5�������������)�Թ�}gnF�!m?հ�����Xl�-�١w.�y��Z����v_��mm���B��������jNY���IԵ]'&]	[��N�?B4��1y��t�=f.˽#b�c��K�m����ϝF#�� ����2P�*t'22f���Eƀ33�K������\ ٟ[��Wn}&�}.bc��C���ԏ�T��5�r�V�'g���HK4�`r�iN���H �n:�4)J��Kh�*[`�g��~c�=�T���S�qc���I�N��ϗ�⮋(Ǯ#*��$������V����k/�i�B�J0��Dn$l֑t�7�z�8�T�/Q����P�ty˔�9R�nw���;Ɏ����3�z�3~�KY�,?�ht�X��Ϸ_��8m��� �I�Tu��'E��ޯ_r�q��e�%^���{����ܶB�3ު�CK�H�+���Ι�#�����H��_��i(����S�PN��E������8T��r=����2�1�=�Y9dA�ϙ�s'��5���D���s`'nL˚f71��Hs�2L䋓'�7��b��A+7C��6�H0�ʵ��pT����k��ll�S�������2ä!s����,���%cD @?XJaV�������T���8��_�lM��C��z	.� ����3�ۍ����F���ī�D���(w�'�d���V�+�]��V{M6��b�^�E���.0��j�Xn03Vq:9Q�-�_�3��`8������9��@�<0$Hc:6�,~o_ D���
�K?6���u��vb�(~܇���t�rq��'�x%���Ov_�x\��,|�B�Թ��f�9]��oUG�e��=�A���|8���a�I��}^���~Ռ����@ɵ�F�#�]蚝�� ����-sG#͉.��`}��@� �;��j��yZz������P����� �N���r�5� a���<
���і_�=k����8[W�/���8�ia��Be,�}+���[�'�����h�ԗ=݉�(���I�����GR5�dg@q��,���I���E�4��:V���5!���Vv��I#��Z�x�r�Wp3���o�CV֨��[����$��oN��Uu�013M~b�����ÎT>�o�C���h���)+R������A4�w,���x@p�W�tzK#��l�Z�tW��4�Ա���Xq-���*
wg3"�H[6k:�2@�0���?
��$���Vf�t�����]"_���o/=R��Gz6G�^jW7����\��}E1D6��X��M�x%r� 뜾��$� �aQHk��\�	�
JX�L�ԟ~]'�|������1��9�ۥ�9;�X'�?�D��Jɡķ�G�%ac���EςwIt̩1�$�XC�^K�r]?[tY/\�k�� ��
�ܞ����lU�Ϲ��2ٿ�Pķ�E�ݖ�<%�����Db���!!Ǣ���v�Kb�j=��>��#�&̃�ҦInǝI�����8���D@d ��nY�9n7�+�DWר� E�M��a���a�������6��?0���t[_l�3L���(����w-/�%�>���/;����g.���%�����1�$b��q��"Rq��e0�'��<A�#�'z�[��Ղ�3�zS4�{y�Aq�}?.
`�o��[d�r2I�p�<P���5�a-��ɑ��5�;y�d�����Ҳ���	Zɔ�>�*�"�-����*��B���B�S�6gϕ^	P�#�	���,l`bS4S��$@����u� �&ͿEJ��� �.&x��0uqD�өT�����<���+�<̨�e��qol|��3�	��9�S�5}2(�@��k��M>s�s�K�s���%�#\q*��CqdY٠^i�Gn��/+<�O����5Z��N��P���wL���x�8WR��Q喹��_���<��ݖL!O�h�0����G.6m�����q�&��f)5Xm:`�f�^4m�m8��(�>H3=u@��߫�����9��~	�P��A�:���ī� R�1ɿ�?�륆os;iyf��� gԆP��e�ןL>Xn�u��� !�gd��}�C�D�0��]�x�p9
�GG�D7��|L��
SVSlTS#\���=��S��3��\>�_��xNR ؞z8`��
������=�*yѐ>I>Vy�ݸv��"��I���%N'����<�)�a���V�����s�!��������S�?Jkh����'qN�w��g���+�A�B�����+�#�5��5��`��;_w�|`a�	7�>��>�WHbˑ��a���~N��R�
�����1>&�����ԇ�������9�w���|Ԥ=?�Z�;e�rޠ�|��οw�$P����	�G17}'��gF�]�w���$a60i?���<Kz��9��nKz��}3�~�az/fO�w�� �+�!�������@��&�UJ @4n�&y�28 ��
�8�AҎqQ�?S��(ٽ(����/��>���`�uf�-��a��P�Ɔǡ �{ S8È.�<��7������{E�D�F��P�(p������u=�3��� ��o�;C��Bƽ�:A�$1�kT��iW@��~h[8T��\���T�[Ea�F�Ռ�<��32��sٸ"��(�6����M\2�w�N4�����J,)lظ ß���oL��ċ���_ȱ���z?�V�5_� �)���z�y'� ����'���N�/z��H���啅.3DZbPX�'�h�u�:�mi�mDmP� '�7%7 S��VB�
J�C��db'9yʾKG�:+�P�@g`�2�Gg��Ht�Z~��a���ƙH4C#I��7�Ԉ� ��:��cqU�q���W=�4�ϑ����l��[����� @�xS��F���||;r_ݦ׭��"��j�Ze}�>$��àd�gW*Kw�}yG#�I�/R? ��X��#�nMQ���*M�md�`H*͖!v��O��vM���DK�M�\�㸜/��9��!?�����\M��89B�2#�ŸZei�(��w��i|�,C)|t��f�X��P+\ZR��0?�|L%��[#�_�tv)
� ��Cy&�]���5�GX|t��7M���V�F��������
DX��vP:����3^�_���:Q9 �����0c�݇�׾ofDfX��>�&5�vo�ٽr�r\�&���_��x]��F}�ٗ���?F50��w�i��K�I�a���<�Y���I?��4���1���V6+2�`��]�̾̅�x)����,�3�3 ?�Ml��n�;d>���hP��0yT�! ���|�'�r����ڡ�Dɢ>\���=��;�O#�0jT�&��xb�
����f4ko]�EiXH&QN)�e|(���&Z1BC,'�!Y_�;��Z�4���y4G����/pD���`�oE���D&���ҡv�g�a��S��C���V�k~Ϳ�|0nt(��:��0���'��"�p�7d�oM9";B��Dm�pZ�4������4�2b��KuT"���Y���V:%<u��b�Hìc&M�<�g-s��I������x������I�a�Nn 姇Z<��X�/O"�1�ee�~9�<�m�S�:e�6�8{����װsqOɏJ"��7��
����jk��n �D���f��?(x>Os�̚f��0��l�)ǹ��|�j��/�Oz {���=��i���pj�@�#��@�b=�A����L��S��r3ǯ4��ƅ4��JaQ�<�_�a�
���!B�L���� �F{�k[���v}rNy%M&���`na�Y�d���,N���9896RV�穎��W�*� �P)ο!��������`������_[���&�U�#TT�NʂWk�|޿�3�G�Ow��b�w��;~L�i�97�7�#���3�s�Ғ�B3�n��b�������> 脦r�ˢǙ�qoLzZF�<=�Oģ��Oo�_�6v���4TJ���u�0������?�1-0�������OđE�9g�9��Z ����
��Aޒ$X���o�j	.39[-WP8>H�Ң�P�݌�ޗB���7�*w\�\����4�N����يY�m��B�/ �/{�b��p�~��.�����v��h�S�u�͢�Xҋ�N���ňLEe;��.R����HGIbu��'�@LKd֣3ѫG��=ʼ��۶l�I�F� cK"ECo��ӹY)���߱����Q[?�5� �p��c���d� �0 �y���7�3��y!qc�ɀ-������%9�s�E
CJ@@%7\n��X"�6�3@�Aw�8�88��)��O������ �E*������93���iY��3��2"|6i��Axh�p�>w8皳�ܰ��W2$�]L�0�m7��Q�96\q�Eʢ!㾳m~���V�\��%�K��8.��լw@/��c�:*Ϊ�P+��K	M��eE�H9!�!��A��d���wc.}����x�Db=������q�w�eM��8�W�.+nw�����#�Y-[�:�����ħ�Η��"�|�M�'B�Q!�|���e�T�]�y��]��i]�����(�Cil��(������c�OI���i�mI�Y2��@V��L�R���wK���Z߸=wzH�9��b�G~^y�\f�O;�e�����u�*ع�b=��;C�,�#k؂�pM�n�� �'�������$���ʉ��۞q�b�P�n��Ж�ox�2{�a�C0�F���f�X+�$��2��}�)�4�!�C�XL8tR��G@1ius����J�M����'(H4���!�m 	'c|��7��y����S�lS"yJr�`>�H;�Zy`;y���J�E��)������@Ѿ�:98�kV��_?�����V����fn"z.�HTfA�*�}���ß+*a���v�V�d`Ca�C�Y�m���SnjM3�,�m��tw��h7����վ�3[��:e����Ի���  �c��~"y����[\(�2*�Mo���{e�&<mM�2s���l��9�����d�����DKQS1���FxE��?�׆�;�����zs�ֈFcG:�{isݱ�?G�$���.QQ�<�� 9)��O�#��ݜ��@,��Dc��V-�E��~E⚞?��H�P[�³��17�$b�|�35c�|��/Q@�Tw�p��#����䎾��?(�����D���Ey���T��h7����Ƙ�RoH��i��3���'��P���G;�����d}�Ea�f^�S[ڽm-I�����v
�ebbxѾ�:?�@}���~tSq���]�͵7�k�yvC�)���L80�X�%fV�s���T.!Z_lQ T�� �pU�US&�p1`�w�S�g���`ѫ�TV�q�6��C��9��;A]N`�D�u�26�������ol����Uh�(\P��Pn�-X���cRk�I�v3��=8&0l�P>��kg���F\�IH�o��y�ǀ�y�����-��*ϩ}f�}.���L|�~� 	_��[�d�C�`˸����~@M%���D����uA0�h�2 ��i)����ЍY���B�zf�m�s<�v����ĆkM%�M��Xz�kdM�_�b
�fQ/�t�N��j������ƇiUX޾��
=�6��G����E�*� ��џ�RR_T/��)��0n�ZF�0�ōVc}��ԭ�u�n��`(qv�����hZ��d�:?=�O��1?��>�Mw�0�?���yb���	<��Jx��0�J/g��3�x� �#�[��C�!�x�X�ǋ����.�g��lW��`����rb;��G��vZ{;��g������|ƒ�x����+3ǃ��L���<M:vaxM|�Q�_�lcv������/T���n(�&���Zd��������F��CN��|%@�e*xp<�Y��{�3�������s��S��d$j�Va�[�-ɿ�4koM���{ �H-?���D��)%x�z$% u��UA�A'�-��Iћ"+��A�Кa92pF�m����u���!�=W�<�t��G�*�PyR<j�]Ì��6]g��2jZvCoE��1ϫn�Aj���[i����n�����V����'A5��T?  ��Fq�{9w|F�_�o��3P��D���y��y��~9L����ۆ������D�W�"�_B��5_EO�W�f��$k3�w��n /��?"�kh��,�?�.�����}�N�<Î��\��/��-	��@�y\S)��Xr'����<��צ�מ~\mk�L����MȡI������#�e����#���z�:3�v�$����b���; ��m�I��! �)������ ���s�`f?L��$�'����k�"���+��_FvI�*[�ϟ�y��غ�Y7���?�ps��j�\� t���u:7h�e�a����:$�؏^�A�c ��+���*!�0⻕ܣs�uc���A3�g#��J�R�p�b��)��Ȝ���⸘/ڍ�7z3Ʋ�"�����WEY��.IC)��s>�:L�,h�&��A��o��KJ\��5�v{9�-}s{�4L�t�9�t�uw���}�r���U���baE+�lM8����.Í�3��`4P�۩=� ���}���ב�T�{��]=t=�+��)��p�o���&P��#�@�v�� �������*���>	�fA{���2��ZW��,Gn)��@N��w�������\Ƈ>"t�Q58����'%y\:ڂ�����	���s��) kw����Ix���+LZYa�����m�6$ͥ�̫�~%�YѲ�i03�T�J�/c��Hs��;�K?if�]�9JS�Iq�Wr|vI$�o?��Vƾ�_�������a�'yQ9��H�y���;/w�*�߇Mb��Y�ǖ�-���a\䣺���H��ϗb��9��=�|����������K]Ag�6<��́�;�}e����F�Zr��+~:������ʌG��瓰����(�r�ݸ����珢�l�V=��N��ڃ5�֤�(5V�Ӿ+�5QW��%4b�G[o���7�|�m��cӽ�~�ِ;���;Ru~q������D��K�1u�ձ���R�h9�m7�1����>K#1�]��o]�-Z�{�kʄ9J'�q�3i���FϤ^��|�Znj�K_�Ώ��a����M�5�ʏ���^����#��&=��M[�7}�U��M��K
��-pi�I+k;���֣�@0��6��э8+i^��[���]r����=V&g��`�*��qLjG�o����O�Pp��zd^�qn�n�.q+�5�!l�P2�=���#;�,��-r�B4*��D$wU��׮��-��S{y+�������wP�LU�i��v�1��:�l�AX<U��'׺w	�E��W$���s�����
@�;���,�w�!d$�l�>�Jp���C;3�Z �|��#~��{��'y��L�;�0�P����:�'y�#����g�-J��}q��XA_�7�Op���J0Z�p1)J��z�i�2u�
Y��ś�j����/j��uh�Y�X��'��R�FR�51�'>��m,#s:��d5��gu�/B��S�Lg�h��@ؾ
������P.�L��h{#y\=�'f9N��.���w&UG' V'
�?��n\5�طӧ������!ϗݓ�N�AR��n��UW�<���o���e��q?�}
 ������y�jB&����Ϧw���|�~^^�*�d����Wq���$�)��+��U��LOB��zk�ٴ���uۖ-���i9K��H��\�����6�
���4<��G܏/L�W3�c���PX�]��e�мOu�=K��-Φ��l �i�xn�O��A҅�l��ѱ���V_�qMK?Wf��TY��?ڎaԶ�M���% �
ȉ�����V����sG�n+����]��F��Nhr:���0�5�քh> .����QG
���:�>��l�[ZS�|���O�,�A+�������R?Q�4\Gꝑ�C�jy���Q;W��� �0��+R6��n�����95��{��򭑀|6�bC4�w�O/E7d����|ïN�r�P&�{{GsT��rMB����&��������5z���\ve���F�@1�yڞ`���f��"?@����<�fr�ϗN�9��㗷���X!�`���4� ǌZ�7��Ѧ�,�I�v���s�	����U	�D����H��T�e��P���a'U�I����׳�3=�i)���0��H�鲛��5���fx��ٗ�@��_��,@���#; SE+��E���	9�'���4�7��w�ɲ���
>����L�e�� ����ͼD7��������x)"�6�d�w��Lj����� �Z�*��{^K>w4!�G�|Eb��Qz��
J�/k���:�`/&���(G��;��8V(?��3oG6���?�-�+Oh#�u�އ�$a��p]as^�y�P3�\� �!�ı�3_��si�%���п���r�]��AꙠ����xv�V=�O�Fp�" �l7kxj�Ũ��h�>���`����y��ў�#���.�֌�c�PQ�>�9h9�ϺC�u*¯œ�L-T��R
n�}"Zc�^���8F���v�V��uos����zj������9��`���kp�i/7h�5pH��ɶa�eȍv�kӱ@�n��ze�0 V���� ��������F^YN*\�3VJO#<R�)js��j�]	Z�����C�bY���ˡ������]L�"���p�lm7Ǎi5��Q�Eڿ�1���m�V��Z�dͺ4f��d��P��4�Je�I�%����P��|3��D��Z�����$�a��Dӵ|�!����ƭ����hwR�F`v�fH6X�;�C9�3��<�y��h��6D���Z� L�k���ZR3�<��_�Ǩ5���\���KH�����a-cĭ�ѫ�"EME����}:��	a�1��[ˈ|�Ty؁�잎n����龧�x,�>x�g��[�ڎ�F:�~
�~�����ܺ�;��xR��mK g���4�n=냉�t�=�v���/h��e�Sr7hskyu����c2!�`6�L#��o�m7������,��2�=,4�}#��"�ؖ��[5��1&��Ih�E*��qGM��N���	�����)bKŌxO͇7�S^z����J�P>L�Z{sF����S5k�V��R=g�6>M޹�؎������ť�w����VT��ߗ�<�u����DQo�2��i7�:�� T��M I!�}>�0�v��zi.b�O!���bؑ���"`��O�q7�'������}	��ۗ5���dK.�h���D#(��� �M�!�<�$�ȅ{�m�����W��N�I�lv�<�ryQ}Ř}�/��Yho2o�<�^����Z��� ���F�w�6��	u����ώ�d���8��~{'����&7�E�����m�uȜ�ZY4��3ܼ�@OU	��ݱ�BE�B[U���_��ϼn-D��֎�_6?�pE��ܓ�a�� />6�(��Y`�2�T�Tϫ��Q��Mbyr˚�����x>G���Җ�߾w'��<�}����#�L�<eH��R��+^9_� f�o͇3���Y/^/&�����[_�}��IM.ƅ�4ț)!LU�s�!���i@�:�Z$X�°~�|7r�C�:9�x��BU���XƟ)v�\,ߓ�5�.�/���QK���A��#��3�K��7�]0
��Lt]�U�BsIr�k�ѺU�#��N%�^bð|�4D.t	19��7��vU4��D �����������6�a�8�t�Z�L�;,wΑ5d����M;��?�Ȁ�0�
��2��9R�/^]��W;�����ֹ
�wR��X��Li�y^�� >�þ��� i��*��l�7��N]�H�r�O�m#�	�^�YV�ē��5����&F��2�� q����.K�Q�����m�w/� {��?����U�M��_��<����*� �2`��������g��ȆŇQ�v~�4�#vF�m��~��X&q����;�:�I㌕+\�ҽ���9f���9�x@~���[�m囄�x��H�j���,H��Ҵz<�{x�s�������&��"��7F6�C�{�7�gS��n9ZX]����*M����܃�a
7�{��*c�80(�nD�ܑ�<��,0g�$��a ¨��Q`��ՑO���7z��*o����G�X���&��[cǙyq|��Z��x�ET��i�.�Hk#���A����^,�IQy��/�N��h��޽�]�73��GV�Q>��ګR&k�}��H���`F���	/�HG����TI���C֏���s��ٺ��������FTAϛg^���D��ees���e��I����a�����٤��a��V%#�n�N�ɧÑ:f��NA��?��fV/���� ��Gc�����@o`K��!h���H@ �ʨ�I�k��I�M���i�o�(�3A~�~��&Z�5����S�6e����Q!s3i��b�������qXXѼJ�~��k �����U���\x��^�klv�N���$P�K�����x")�g�v|{�z{A8t���Lz����b��P�3$/$�����翆���j���	��z�)0y�*��j=��p{o.u�c6T�"���#.\]3;���@B�������v�-��op�%�e@vJ�$H��{}rvg��WE�x�%�V��&ai{��`
����+���S�F��ꓚ��p�[�-��}�2@�������8S��cAY��m�(~�;�g���{��!�k:31�C�4!�|P��L�kF��́$�h��r:��y���%�����x�)
E'�"��!:&_�i��gy�% pF�k)�l�H'�C`:jҋW�P�S�O 3�#��	~1��󤛴;�i�>\��C�$�`/�-������n�L_�e��ӻ��1�{��[=��t��Ô����<Jko�O��av{e\���NF���-8�4|>�u"�+����V͛b��������S��0}}������eN,l��ī[6�4���I�D����� 8 �������~N���5x�R�D���R
=�el�#dM),�;��:zo$�A����i��P�<s�n�ؘ��x�"�}3�撁�(N�h�e>��b�cv�S_�|*K����:�����T~S=�s���M+�6:萂�+Ʒ� _ׅ�̥�Q,7�X��f���s�"F�gh1���ч?Stf+f�_;��CJ΅0;��|�}>̀��+� Ġ���#[�=�uQ��R���RG��ֹ2��Z��&S����QHf����w�Js���f��y#�~u3b���<�|�m��>(�rd���=P�T訰%��|�9<�!�p�i�_���c��13;�l��Hq����[�<6p���c�5���/�=���ָ�懪"�|��kMfoc+1I��z��2����g}o����⥰�Wn[sW���O���Bʕ�ۘ1��n�)nMu�i�cK�r?��[�Q�,k��&TD̎G�^�5�^$�\xL�b��+(R,
�MH�G	'��<�^����s���O�noA/uB�8#���V��B_J��#�hD�zM�[@�hL_w���^�$6hj�n�Ѧ��ҏz{Ŵ���=��F�2_���Z֔gUC�o�2�� �)�*��'4�^�$]tn�`p����(�~�֏W�KZw{#oڹ>�}G¡�,ϕ,���k��.��q]4PZ�}���xsLL�+�F��2�iM��E�]�&K�e�h�c��ǑV-z�x�
jgiZ�Y��N{���{a�t ���O�V?�po�O��&N��'��K�K�������L[n���9c��fRXH�ɛYmyd!o�U���j4SI�S�U���
��N4�c����Z�̈�^��Ұ����F�0��p�|Nķ2�^����m(��ALkD��!�L���$��k.���-Ey6����a�3��>��Uc­���9bВƹQ&������N���F��0W�Gu6>����{u��j���Rk6&��^~�@��5��D� ��KO�T�u�u�G��R������n�֬��u�@��h�}�(��v!��F�u��a�l'~��2B;u���y� ͉�cO����n4,�r{�a����ͼ�cʕke��.���} �� s�y��z*�b�ǨX�)���ڐc0)���O{�8�v�^(�vk�Ā�Ll�ꦗ���`AՋ�س<�ǫl	a�D,kr�VZ��
�jt�&L�k�,�酿��4�/��}g&����ȯy�y��$d<��N�67�&@9�y�u+���U��n�k�<O<�r>h����6���vۨ��5�j�^�/ئ"��,ԭl�/���y�<�
��:�d���A�r�c�rM$��@��a�L@x�[�YO��Y/	ol�w
rZ�狩��r;P�G���|Jv�&�.D����9XX�?���C}dS���ڶ;�Z�����: �"H��b�,��}ڞ�HQ^Hz���$��0�
"~&�ǆֲ���h�撋I!�4����Ͳڏ'#.�c�7���ס�	�}�t�>{E%��s�Sx�:���
���@�����B�VJ�����4����Xr ��W���<
��^���fU�t{���o!�H�#�>3}�f�%�����*�E�/?�1�Ez�ůa{�Ïe2 >�5��� {�����#Uu�U���y,Ϧ����m
@���x��'�6�@��8:��8���4!#�79�'��m���"�s׿t\�ⱛ�5���\ �g -���:�Po1���g�pA�&���'��+Aާ>bb��).�b�yB]n�K5W�\El������򗺪OZG�հ0a1�<��,6U��h��&m��w��S�J!�m� QZfVO��z��z�'�z� ��W��*/�1p:w��l��@���%޶���/�{�v����[ǜ�����T`����E�G�J����0�Ԅ�N\���2�_Kh��-?:�8VQ����.�z|�s��L��.�t��P_�f��vBB~��P���e2��w�:����.R��R,2���H�i1gY��^��-ȗ�����nϽ{?�����������k^��sI���U�Sӆd�eq�^��Ro]o�-�_��>�����L��O��y��Y��%S��48�|���|�<[��韗F���[>jǙnlӮ���b����Lhَc�t3�U�sQ�j$n�љD� "kS���˥��$eA��ٺ��*%�Ld���*�H|P�}�5[�7�\�O���	r���[��^��~�a� ���Vb�}�@�nzV[��"�?�"�∜���&vܵ�6�m�n7��t�����rl�bA��w=d'Df�k��7�H�pq"Ւ䛫���
�J8Wy��E���\��FvI*��͹�R;5���k:^� �P&x��� �����1֬b���H�w����~��o '�7�����|O�3��L�x�����o���AG���$̥��K��>� �Ջ��@P�yA����/ו�\�d9��8.��9�f�ణ������4���^R����*�ʂ����%ִ̑jË������,.{)�/[Jv���n&�'P�42}��ZN�ZUָ�tzET89q�xFȍ@�5�Ȳ���v�@�hd�V�^~�����a��?^L'���WUsxg48�Z�ַ3Wl��y�� :���Lw�,���?�{G�&~䁴��M�����,��O��4[4�a�/@�2#��tK��C��΢�a�7�aa���Z�^	�4�"l�����G�YF��5[ww��.�ݝ��$8���]�Cp�`���=��s��[�_�Y�f��T�~v�陙��O,�Yt�=��)',�ط	�)%Ca����ͺǕ���8ܜ�Mj�R9m5s���_��h�~����-��m�yV�D�;���?���`����Ay�)����t�$�[�m|'���}����/���J��5��0�٥�x����dܯD�z�
:�O���̟�:}���}��XL%����dސ����q8���/� �?�c%�U��	���cH�X٫yE���#�Ͻj��O��K�#�GV�'��J�.%2Bu�W�E6YD#�"R`�r��h�gOFV�c��C
�6H��|J��N�[�+����� �v���C��D3nsyuc���^6�3z�7T�|���r#B��	�=
Fp`3E �H��Lc'f��d�h������H�+�H��p~���ܺ�6��z�T�I_({T�p�+W���;s&6u��.����aC����o�CWx�+��(��0PP/=@�n�yo:�n�}�|��[E��S��R,R��m�	��g|@��t&��ͧM7>'D� J����f�tj09���sf��Y�Y��m�ќ�����>��w�����R��@	]�=�컽���J�&2��Ŏ�� ����V�����
?:_��h��L9��QxC֠���9s�3u�������Ì#E�*b����@3�3��aˍ��E8T=w��Qa??����`=h��ʛ_g�̈a})�)x�D�<z�`��ӝ�y�	��n�ϳk�n�&錓Q?��Ԥ�B�  =��:bI�b��9R߲�����d�5ڻ��/��]m~�?��:�2~�r�֓�Gӵ���LHW��T�]_�L�pwr4矙���'n+�wogqn�Gd�MQ�#�B��N]B�4��gp7Zw]��0��<���A!��;Z��=�λe�}��˛����m+@/.8�Ƨ�����Z�b�&e�>q~
��ҭ���OW��4��,��?�RW=Ԇ��gtA1#�-#ێq�q�IC� ���d�b�.���1ccR���$������2r���뗞򧑽��(�-%"�\Mk�,۱����	Rܩ���$P�hk���7F	�0k��#c�ՠ0�@��^L��X>�[8<�8'�컊�d�A��0�2à����p��#wU�@��E���`�#��\h0�=8�n�!�"��8(F��Ť�Y�p������X�<'�T�JT4�$Kn�>_�(=��wO�3�Cۛ�֒�^5۴�M�Q��Ъ��92k � >ɠ�D���9�?wI�����$��'-���1糠��N�S��3����K�v�&4k�X�R�T/؜�7hPb�8N�콃����*8�d}�P�Q᮶ �U^�|����ޚvɩw�E��K��ov	��Ʌ��`X��aX�S���+��>Y�8����,�O�o�B%��l'���8��������Q�=�n�_�m�eNڛ���͆���f�3o��$��⦌��8�7OMDB���7%�bz���x���]m^)��Q��<�q��A&�B�f����	
S�q�?Hf�G��I�3 � ��1b��9����s:���;�
��u�X$@aeb���2[	$*@�3x�S�O唇��h��1�{fd�����
.�'��G�n9%Ss�Ê��� 2Wu�B�䘏��/��caUt#���U����.���f�Ŀ9mҎn_�Rě1�b�u�t�C��N�fcF+w�[z��I�^��,|X!s��Ɯd��9:�7&ݯg���c���o�j�����R6˼I�r?�ɨ&-)�i��ęۂ�x>�(�,zz\�����0���	tۓ6��c�&y4ޯ�Җ�^,�D�?�"��X$L�F���v�,�P�Bo�7��Z$���P&%t���J	t��T?������|���a`wo� 1��3����MMB|�>�������(?Ƅ�AӇ��7��?�~���\��*�SK����>��X��˥�}���g$ui�����+�h��D�{���ccd��p�i�O�8��|�D�.��x�~�.⇲&�W��k�7��{eS���%�a8|_��3��������'��	, ��ԭ��5�dչQ6���G9�$�8��`�A'��W�w[�Jp����c��ϣ�_r:�E��$Y�_kLN{�J��"��Q^L��z��V� ��nN����CCȿ���;d��k�/�T&O|��k��h��E���m&�V<����ݻ���;g�!@3���dQE`<p����aR�?*�e���W�@�	���?���y�868�i()_>�m1Y��r�?�O�O\T��6tfStm�Q�����1UЭ�X��8��/�GB���撖��������Z2��:���ſ��[GƦ�"�e�	~.3��@B�_�߅$�gW��=vs�d�}������.k�Q�V<�h��k�w&b-p�3��N�"�f��%{�вV?���4T(��|�c�a�����X�����U7�G �Pj'��Ll�q����D���������K����$k�(�gh}��3��%:�3��zӚ��ր���m�F���xy�]�p^��Mu�{,��ͤFˇ�QP�����2��{�ѧ,lŌޛ�dĮ��8w�iC����/�Gc��&4Z���,��ˢ's����*EBEN]?)��� ��'e�R3o�oT�bc�	OͶ-*(^��ƿ��ȧ{��{1�΁��+~���`��
Y����F������[��i~��d�!y��f��_h *r<��� ��7mg�S�@@�G֦�nr�b��������� ��v���|�|��;#Lzq=+�眡'�CPI[Ԡ��3�i�V
�J�_h%P#�g�c��OT&0)���~��8��%yp�l� 8�J���D��$uZY"��j���e����r��u����"C�?'^�*��_}C]ͧ�`
������ � f�[���	����a@����+�r�	n9W�6[>e��*�w�τI-}�̄v����l���7	Rj�p�i�bEX#T�4���a��!����H=H�V��31Zc�=���b�������8t_���B�%��Zaj}��lb���!{B�IF`R.��dhH�Y]e�jH0��.o�t}M�+��BS�yi�����j_�1�B�*3eR�l����E{�j����J����E�dV:o$��sO��ы�C��uy�Tm�ɩز�B�C�h
���r";)ь�Q��͟��V��l�w�<���F��$H�l���9�H���i��S��πL�p��ԫղ��pG�����F�f�P1sg`���G��d���E�nl��S�M@�a3B�g��_�O�6T#�'<v����R{}�ac��{,�r�	$r�둈S/�3� ��a@�3Ki��Az)�~'�� �G�TUF?g��uy�8�*o��D-�����Z|�uT��|���K-�l�����c�P���JgǖğT������m$��n-�Wqd���2$�l⻋����R�j�Z	�;]�S���Pe�fϵ�� Q��6|���0<ot����3��;g$嗫�����%-��t18bв��,L�|Cx�p�Җ%�QϘ��,�j<s��C0A�V����
c��t/}��ӣ�8�� �x�������zc�3X+��!Z�a�|]�ކ0z/�N�)wh�ﺧ���q��چ�u`訧E�?�;��u��>��AFV~\��a�L�i&�S���f���|��f}�7K����ˣX�{A�v�3��q&�]��Gq�~A�taذ+آ*V��9��h��A����5� ZV�]�r��_�;;�`�2d���RqJzpc
���d��������kr>nƔ���w�7T�QԸ3ӇT%ɂ+h��@rvMn���LKsJ�c���ݣ����ᒼ���H4KN`gL~G5���5ǻ�u%cz��Ι���u����ͅ�
9��6J�_�S�[!'����qx�i���8ڻ����{����B���DDL1&�Nx�fv�Bt��n�d4�C�Q��Cwux~`��b�m�BV6��9	���(Q��sq�{u-��w�Z�}q~�g�<P>
��2��Tc��^��g2��P�69Y�И�.�E��o �#�0���R��R� �Kbk�@	Q�y��nz�Xo�T������YK�o�۴@&�͌`!�%MC�鰥l���S�W"aJ��E��n���iՖ��6sƋ}�AGv��#�
	FPq	;"pZ}a��[/��c��"�V?���eC%ؗ�<*�����PG���OsSNM�Cq#�����O�7�>R�p=3@��t��x���[�6�
��
�Q�2����s[�Yi���t��Y'o5�p2ryM
�q��Y��Q,�@�161L��6��:�trx�Qç�1�6[o�l���8$���9�"qd��"Pkr���]\y�IV�ʅ�u]Q(�#��ͫ���� z9gV!�/�D)��9|�4 �'��⳩�_K�k�������~�����~�B�{?�v��8#0EsӞ^:�t���!_� ��<Ls<Q�!�0��:J���K���ӧ$tS֞ �D���k���1��v��,���`���M��r+�A�X��n	���^�gkcV��R��ގ~�U��J
�u�JU��D�_ޗ�;\Y1�M��vQ7�ޙo�vm�;漿z��>��~��+;���D�݌��W��얗��Ө���ўy�?6�܌��,`�����.����jN��!��>8+T_�gK� �	oޏ�����^#�Rj��%@��N��W������j��D�=��*���c�6j�f~�P��`�6�Іk�rϞ���6:�-��[	���G�����">&� ~:e.�j�� �F�5r/d�E�����}��ZH�3h�[��<3�� �-��d9�6G�o3\�} ��m��K*yb�Po�CT�Ԗ �J��\'�XI,%�]U:$u���4�2�bqS�&3�k�����Z���^�����8����y��\���L�3��*��W����#�:���IBw|d�{��
�/�1Br�]QCrH��9��y��
O�L?��ôa7�fc4΄��>��r������G&{u�︐��r1/��0��$��{5�B��9`A����W#78ma%9�ו�}�3�qrv(8�{{�WI��G��ֆm-M��ƹ��;�����d���l����nR�D�<�5�5�0Z�A*/ԅʿ��:R��D�7��ՅC��$�*Yo����E�
�B���}��$Ml�R+�w��# ��$0g[!��ɚ�P�a�����EBº(QH��Xl0aMD9]�	Hۃ�Q_�	L� ���Tv��EhY��C�,������p������ �F&B���Y9L�̬檘UՕSy���;��:a�I�Gx�+��zs����؁�E^=cW1�@=��'�W�v�{��q�ο�LD�ľ����}�⦛]z�t�/�PЗ�y��$"���1�O? �f��ް��W��/0w"�5bGR��k���@����������@�p4�l��iꢚ �f�I���*e�9�z�*�Sב�	��<a�&��	��E�����`P;�}��|J!
�L�Ά���jީ��aف�b�ϵ��p��-i��:�䥱�z۫�2bk8b��o�IV�sD��n��qp3�pT�9��%O�`;:ڽ\��n�
Aݜ�����Y��/hdz��&�݌�e����~�Ri����d�e�I��٬a �<ϷH�Ǫ8�t���j���S`7�E���I6ԲoE������0*7cS#�J��~�	ꤰ��^�x* |2!�Y�iڞ��<�����1��p�Z�B�|*q(�?ӊ<�\��&�E�up�:�PAɈ��M�r�����.�y|�PܥR�s}��+�D�1NY6"���
I������n��s��+�N�
o�g��²D�	[�V��EdN���z����e%!��@�Ó����0?sJw��2���ף9�����`�O_p<�[�����-�cM%W�N'^�G�����Pf��>S�lbA�}�]�^�G���I'%�9�
���m�j���>\��dFVo�Z,FC�����-"K�h��.|��|	zD�ן_���"0���Ő7�dZT����1����~U��ax�z{*�Z����튮�
�x8�F�\�����,�> d�吇���Kh7W��
W������C�5����\���ON�/�:+�gq�}M��^�AĞn��Z�~�\_'�d�*�h��F��'r7�Ȥ~��LGp�z|ɯ@DPs���(��0�L�X��i���e#�)�c:�.���ՃNz�`&=J��[��R�s�ۅ��`)^L�/r�a�u����T��@P~5�H'LFV��#��$�`�!3� ��v��xw�")OV"݄�;E�r�W=0�ϵ�(|�nc&a�t8�ߔ���3�6&�|I������M�.�fL��b��fk	��/�-�������ja<���4��TV:$�����m��}{�"	�"Y�8����o��A�Od��@�~���^��w��_S��^��t�����1H���F�3֡U,���ɥ%�ҏ�M�h·���n>{%�ƴ@A��t�ۛg�/�˭��C�����]V�ڡ���j�CgG�U�Z�*�M
�>Bt�n�[��S�
�f2g	�Km����ODI��A�@u�N���옿TM�s�[v��d:(jI�+��\o�T��۵Z�rt
;�ɷ����E?�Ԋ���<�����;g��V�AqY�V�}tKH Cmd��*�V��e�F3������ `����мÐ�A�D��o�I%�ijp@�r_ȋ.���M���ޮ��<q�1��4F��۱||����gJ�õ�A���#��/'���}p쫢Q��h�<��Q]nc1����c�d�	)����ڵ!?̃����'<d�~Q8�'�6��ܛWp���\��c@"���׏�t �c,����KϿ#�m&ׯ1�z��e8t��P����%�����޲��r��srܛ�"�ڣr[6.[1�+��`�GЕ��X�����	;����fEd��W�銒��x/<r;9m<�k�z�K��S����u=jyJE&K�(���67���6˺}Z��7��S$\=o�n'����M����UЃސ]�řVeݔ<��W��8Myq#���ՊH������5�vɋ�o�	X<b�x�ުji�q���0�ef&���gB۱���;�$�����ӄdy�-a�d}��!���jAI��b٨�������5�K�K��`PLQhr�5,��utz����>�0����`�I����	�Y�K%K{ف�Ǔ�������d�57��;t����(X���$܆�}�3/g��!�F|���#о�T�@s3�5� �d���)�)���)�w�&�)vdE_�f��^L�ZH0ȯ�޸�m�ϪD������wU;��� ������#Хb�:.v�)�<Ŗ�tP;���Q@jҩ/׆Qrg�b%J�%<�W/]-N�t��B��d|�G����MWzq�2�'�(�˄����޳>z���R����}�ٗ��"m�"*����1Ȑ񊞹�p%;��-Acd���(Օ�����5����d1h����z��
�&x�F[�Hu�u�%Đ�܆̞�l�x��~�XK�kL]~�4em=��D[RM�M>�)��椡<Y߶O�F��E�N]x�*�w�OYeGw�u��j�h�xn�M�_�w+c�\t�~�G�9^����}�]DSJ{�~%q�Pa 	I���p/�>I�kXd7`�������|w�%c;8�4������[ʟ��2��ݦN3">�j�QE����L1����3`/ng����#Jk 57�!vT�!i�2���7�l��w��ȣ���ׯ@c�aQ�f�|�2)�KY�Nv�M�@VEJ��U[�hMt��C�ڣ[J6�v�o�.��4w���p�7O ��!���:ǖ"\I,��	����3�f�EԢ� ��;#�)��8��! �>�/>�.��2Y�ߨ(y/�P9����"�J
�02BNv��M��냶p�����)�W�c�Ǔ��ఇH{m7��x#_��̨|5�{�[�;r����q�gg�L#l�ڷ�Ț���v����N�*�O@�)td���b�l"�z��cH�ɹ�5T�圝���6 �g� ����"$Q�h���鼍������Υd(���Io�B!{ғo�4d��Z0�d]�,l�05]�-����� �C��L�c�^!K �C]�Z���l��i��Z3!�9�dCW�R�xJ�5S��%�&�?���Ѯ�w��ᔷ�G�a��������A+	��K5��فl�,�-%kR�����p}lz�:
�D�]�3<V��+z}:gC���5�e�á��żǽ�5Ej�4����>W���)v6�G�A5��B�j�E,��>���U�n�-�%��e�sN6C�e3#n�#��dhf�� ���1���{Z�����[Gi���s��k
����{F�<n
�,ֶ�$-ωۤQR~�F{P���í�R�ŘX�_���Ҋ~�̽U�RCN��7��*K;f]��J�����I�	��0fhi.��j�IV/dP�|g�i��	��M֭wo���u?Wu�`%�*^j�$ȩ:ʕ�'�3F��q�%��E�ցk�;6�)�$�b'd쑚��l�F�`f!v�_�ڒ7sOǡ�z%�a�SuO�]#�ˑ�����xj0�(I��$�zF��o|�?��܇����tU��.V�|�n���������^��5y��گf�v@]�{z�rv�^!B���N�(ؽ�=�<
�����,���\��T���`�SU^Mܠ��헴�a8���~d5��q��ֽ�,)��v^��~�p�'�}öЛ��'�w���z�zg��yr+�CYO-&M��F;~�=�2ߑD!d���/��/�rP�c� �9 �G��B�4Fg�N��$/D�Xd�Т{�~I�H��ܚ4���0�������|h�֒:���;��:���y^w���c5�ce�LC���Rk�Z��ο�O�E,�yN�v^����2z���+�G(X!<��,�o���,�u(���3VAh�>� ����/��f���؃��_�c}Dz���FP2қp�S�I}:2�n�s{x;��9�l9RpZ��� ,)>P�_�\��d7��>'K��ߤ��|{9�FDNW&�I���-r�A�*���ܮ��]Ǯ�
��ĵ����KM��eܴ��։�y��Dދ�K�������3�4�Ҥg�f�̊I����!���]9GN����"]�[��I�������/|���5�7P#t��J����5��RV�:�⎘�}C�����.7n(~[��n�&��ٱ��;�,��Y�Ε��������t�M�,��:����%��^j
W!��K��@�Yb��+~�,w��BV��7��\N��-b�Y�1�HI�(e|�d���PN/�����%���=i-@�Ԯ�,Y�����ˉxp�/|~z�<��$�Z#�>&qr���h����\��4oc* ��k�`	T_D���Gd1϶_�ŋ֎��!DG'��E/��1�O�HT�t�L�q�o��A�O�~�u٠��Rz�L��*Zx;�G�����l2�+Oz�����	`�h�m/�(��=��7�RGe��ě����sr�4WlC� ��x
����ɩ������@C?w���*�s���W/�#�����.�	x���KaK�L�t��|l���u��`%)��0H�V�v���
rE9����C�T8qZ���-Ґ�'��gE�@���;�9�qR�I��1����-�K�	ބ�&�����d��|���O���H�Z�V�b׃*��K�r8�I��9�) |h�+���+s�nw����^L�^ٔB)o�$�E��1��\���%ƃ��ƙ;�?�6>�;�/}I�	c��Hv攀rIF��!���m�������겵�5
��w"k�@KT-�Lc�35t2���4�/3���6��[W��>K�l��C3�����ƫ;�-� ��0�������D�9��5��0ڭγ��"�]`��c��X�,9��.��n6t�~u/� 0Ʈ�g����%.\����_K�t����u	=%�Y�,��h;��6I�������^$.�&�{�B7�����뫳V@gI>tg���ұ&)C:_o�&C_ٌ��q�߈�������K�q��۔,�ڦEa,F��� �d+��Hd���-G��!i?|m��g��֣sb;dǵ/ݮ�}�H��3�vF��7��Z��>n��$��J�Y�'�UR���t�f��8Ӑ�`����߁�(�ܗ�`�����Wn$Z�y�V\Gv�
®ίڻ&�zv�v��f�V�jT�>6;=�殠n�2���Q����Q6H��!��:���
���/8ST���~�LB����>����Ѝ�έ�����|X���k'u�����`96 <���t����\����P��kӋ��e����1K�V�"	�I���<׬���a!5�=Z�q������z�bؾ����昵M,Jܫ������O�-�t��\���*�S^ɲ�-��jh��{ٸ��s�p=�ۭ��'n�mn����v��o�>��D/��F�����U۴��y#�b#��1���v�|��a7�@CS�/�s�-��Ի�d�1ߓ��� �MX;�!��5���^Q�f���1���g(l0M"�5���h!a�������T��_���̖���zJ\Ga�؜�c��vܐYm�Jd���񴼲œ�䧶'�C����I�g��ē�\�I�j�ؿS�f�vb*��3�i;���V�qʔK�y��e;�=�I��D9"A�m�Is��z���ޏ�
�1ɼ�i0؎Ő�:��K�s��7�ن�vB3js�$�'�n%�3|#7�_�b�&뫣��^n�]�L-�Jt(�3�q���D�N�������vN��j_>v�<.�*��O�.
m
�����tu�aE���C�5��]hI��mR2%�~O��+�f����^;e�����d�}	X3=J��>�@4��?��O���U}}�X�s`~��K¶Y�r5���@@��H����u�����V��_G֧����\�2"�HD�5�g_QB�Cyu}@P���T��wf��%a�~&��<�B ������.�����5�S����mN)���D:6�^s�r����B��H��}I۸+L��K®FR~�N��9�d�cxמ�Bn���![�ʀ,�\���*���ߵ��/�|��A�� <��y�@ǫׁ
ג}���<����ӝ2T�~���_�`��GH�6!�n4|��.�D��L�k���epQݹEP�����mx�r*��D�w�Y��o���t�J�^4��S�GK�lQ(iE.a�M�=5zi���w��	��"_����i%#c�sC����j�M��1_o�|?g�w�l�N�5C�K�36_�=,�2��]�&�y���Ďl���z.�P�	O�jWϸ��(���I����2 �Z�h�Žř5����@�$�}�k�m�]�X7�3��"#E�BOQ�r`�� ����i�� ;f(5�����3����_H�c>�K�\�|��������,$=��]G<�M� �oOy��P9�j9.k�_�]'��&�R|�}�T������oDH���XT���a��E� Hs�d�6��$.[�h�T�i݉��z.��%Ug �������:ۚpWF�r���fz�I�����f����g7�6k�����턾�zQ��*Q���i!5#�a�)p��C��bo�ݔq�����@�m(i�z��[��RHܜ�bc�������&��&4��>�Q�ѱ�^��Ӊ�>�� �M�A�5��(�ym]
5'8O[���jG��l�s����y��8}�x�ʒ�����EM���`�Rg��r�%�2B S^�7G9 ס*�>o���h;�<�mT�Y�9H�J�a�����M+�(�T���l����A�"��9���x��j� 8I�WX!*��r�.хl\7;�o�+����N�Ѯ� ��ـ�*p�@�(�6�UG4%��A?ܶ�����׼Y ���HȄ	x�M�RV���mJ��& �X�R��J\��?��wR}Q����a��	HI�W{QB�l�ُ��Y����{�Q�bm��r����N����9b�lɺ�8Klb�>�*���H  �����8��.t0'��bg_�p9��㩢*n�����un��WݚT���k��jΆ������K�d��T��Q�.Y*�����{Q����Y�tY��īH�m��M�[�:�@�M�(Iș����]�"xP��m��o涶�{Tt�x����<V�F?�#@����{�
Ŵ��^v�4��h��U��\��Ӯ��Ż�D;�����95s�}yHW��������V*�NEpI�~��sI�D:v��$��	�0�/۱7D?�^B؎�f^�U/�q�Ѵ�����.�Z�۟yy~��3�P�[( ����j�O���Ҟ ����!� ���Բ����,'���	C���"�
9��y�>��N=<l��W�1���2����M`���X�U��xJ�&1j"2'�����`�K5�:uB1��Pʤ����ިr�P�1A�V�Y:�_��͘0�$���P��;$�B~���s�-牖� C�Y�m�G�f����b����J�MF�� �R��':LH�L��}��	T�M�fb���
B*�/�;)�uBk�f���Y� ����FP��^׿�ϥ�0�D����%����?�X�:�4N�0]��#ks�3�����ц�=��n\��d7��A�#���/��\���s|�Y.x�~��̀�3~;ߑ��8qW�U-V���Q
ȟ08R�lVbߕ�:���y��U�eGP�b��?ږ@�6k���t6{O^"��B�x`d�.ݽ��M�xw�k,|jj
1@��9V|��;�i���u%����bi�b"=�x^�^j����"	ۈ�0_$U��]������+R�k��ˑ6�z~��c�(��I:s�����t�5nPX`��4m��<�j�1�� �3���=�Z7$ԕ?�c#�y����q���I8�{�kxmė�b�M���7�6��,uOK�����j����剩�u�C���O�*&8��4SC�Um�yu.p��T6<����d���0�0��X6�H"�q�7�ϮFDx
��)�^�5�0��?[4=^A�?�
�X��5zٜD ѽH�찚����`�o�~#)��L?HNn��I��*Q�L�n�5��&
�ۈZ��ٷa)���K�/�dG��9����.�fh~S�R:�b]*Y1%CO�e�F©��	$�>(-��.�Ɵ$����=���E(R]�0{0~������&��.Xp��vO�б=%���!��b��
�cz.3n�TU$j�?���׊j��`�ī�`;�ʯؼVW�ي�*U"-�0,yaW�� K_f�ސWWN���Xzj%��(�p�E�a���C��u-�t�˗��o+�Y}�+�(�q�Ic/�lP�t�q�3�urL=� )n�
;.ǀ�3���ˁ�C��µ���&��
�_���|��d�@^,���s� \���#E;��ۧ����;�0)��/{���I�>��`�jՎe7�ڻ}�ާ����8�x��T�ɴ�N��5`۳�^��d^�O��'���O���/A�����/�j������%�0����@��!!�A3� �������C[tZ�I�OmD)@����oeQ����P��VSFHQ��{�6�A^
�<D��Y7"��es`�J�ř���V,��������?����U���m�,��O�ίV���u�~<��">�dz\~���]g����TG�l��(�����~��:�p����\`�#�͟\�����AI����:)����47�R�7%U
����زc�̸�ڨݐͷ!�!�,ם�ۣ#��2Y4M4��ж��gmn �v���5��_ޜ	fց��Źhd-��[��W�{�Ku�hn�^x��Y�A.�U������]���I~�ƭ��������������"���ܝ��J�)2%�AZ�e�5[j��Gx�ΡڇD�GD��p'j�s"��}� �������6s^P� �r��@�Ҁt�ф�3؟�`:_ŀ�d�QZE�2��S(�{n��h��>���q�	:���P�'(��^���z̵�.7�:?2��������}`yv�G|�Q����ZH�,�W١W�؜�1����I�>�_Ļ6gCW��� "u��@E��Z�n�~�z�v�5�T�����}s����f��;��M��WpSh*2�/�Z������?m8u
���0|M�5�,/��I��V��A�g����=�,�.�:��O4k�ja3d)�]Y����0F&���#9�,��z¾�<h�3N��A���Q�`���/��$kx���_�t�SG����:R8
t�ڏ}S�meЀ��^#��ZmY���md�?��p�2_t9󾉶;r';Up8��8<��24H[�����z��A���E�:��>����
��]]K�RvQ�%���&�ѧX�a�8{9p+^zZ%�զCs�s|�����^!���e�v%�~o�T,�!2TL���U=����|�w�Y�nR�\�)��Frh�J�2?��ࡑ����#2�M���Ѷ��}��즻��0$aW�� 6Xc3�rtI�X���y������������%��Ǌ&2n�~�,8�� *ޜk�B��후��s���3�n�LL�̽U��=�ZZ���J����\CD���z ��l�q��R��Ǔou��s��W�eڹ�F�b4���y����`�{7�#q2����#O�^pa�dQ��r�nQ*�3T��
�a�%�8)2�q݊�c��Hhxr~�脷��ُ��j��f�!X�:��]�n�RГ��(���>r,c�-J�@1�o���B�0V]�P(U1���h"�H4-��{m\(�'���P6@`I�	B��L��@�`,2=ek
3��ܾ�=�)�e�jZ�� ���z�	���|���� 	,��I�Uq�f���L�ܩ�bi�I�2�X���ufژt���*�P횯V��K����sǙn�W���� q�	���p�
��	����W���Q����(���%���cKy�?qy��-B���'�йs�<M�t��6��˪��^��o��~��'�l�"P r�n��,*~�G)��v��m\z��n���YH�g�t1���1�e#�}qE��E`�5����9�b_�x*�^���X3��q`F͒�(Je0��^~u ^6ä��m�CQ� ˻����-�����H��ϧ9'��/�@CdEA
Q�0@��ЄlqŦA�@�A���t�B ���Ѐ���+#���twb��r$����Hpn{�E��w��������k�' "zM��h@���n�dz�%D���ey"�p"PK�����Ɖ��{(��R���K��@j��sښ���<�Mo�L����h|���e 28Kqh+��:6�V
�ʖ��YVj�2�	�[ٗ�rr
4kZ{�A��7�����y�콽�C 2M7�=�8�b]7;���V�ʅ�%��P����Kg��9/�XT��"\�m�-Y�]Q�W�mu7ε�J'�0��e�	�YƙF���җ�n6!�[]y��U%��0Q��7I?dWo�#���v3�T�,wK��ش���T����1�c0�uV��<���n��kZiC+T�dG�v�#�TFWG���&H;L���*J��R�e��ppCt?c�!h��W��ɗ1Cf����(X��@�uY㊙�5�MY���5��={i|>���e*Q�Q;n���F_�立%2�~������U�%���H�E���i�5|�?p��9��K�K�ߔ����0j�x>��p�b�BQ9�c��3����u�I����2��Ks��hŇ!*����W���1D��U�)b ���),��o�r���XZ�5^�Y�SL:����<Z�����-2n�*%q��jw��Ĉ;��s�2z���Kiܡ/����֧��pB��(����gD2�l�w�k�q�����F9E�jE�B�tʿ��*��[��#�ƛ�X�f�%MV��ɶ����P�
M�I`\:�.2o�����	��'٦.9�<�u6&\<��#���� �N���l�o��4��á����E�Yi҈��F�i��,�,Y]�>׆n�ςgF7Nr�Ԝѿ-��di'�<��U>�)^�B��ʞA(L�rȮg�p�AGYKlCS� �����տ�׼h���N�f����Yj�N�篲K��8 �S�݆0c�悢���K�?I����t[V/68{.X��K�/ۢ����|8ސ�e��Y�dQ�%w�<�1{f�k��=c�ѵ��nF��n�z꙳R�?�]yO{�T=D J���H" H�m{�����l� ����-â�ڶ�ABA�A��n����A���n���$�a��a��=���~�����xg��X�8�c?�}�k��R�퍣�rľu��t����U�0�
��{~L)�e�Au��C�ő^�j�?Le��
��e�l�����5�������%�w���U������=^��)���>��_�¶Cnr��G�D%Kq�f�09�����C��r4�C�l���a��ɏ�@��|]X�����)��Y�����m�`���47��5�I���}W!*#�߄�׾�P/��i��b�����	�O���g�4U.wv�l2��Q��NRx����cA��[�X�d�mq��ZlE�!3� $�x��@�:
L�*.�g�������X�&ʷt�Uu"�cj����e�蜅����p5����>����'9��J��*��.�"���{%�+!T����o�>��2[�Oz!��&{���|1�j��2��V� �~�LQ� �П�@r*�������^��h2�W� $#!�~�9E�]��'�$Z��M����J��&eJ��P���Jd�\[�ƨ-r��_-S���@�-[X���w5%��0�����53c��aW<�M�� ����kٲ�ˣ�y��P�Oľ�pW:��n�P֊����7	�A����(|OR��1ЌWW��W���]WVu%zm�n�n^t�i۝�O��gd��H��V�r�vą���I�F�&��X?��Vjf/(?�!�9_���x��g�=q̜�<v1�JԿ���ӭ�&�R����WSz`��J�<,�ӫ{R�.
p���;�H�S��e��cu�!\��#E�	�%^3`���k�唥T�	ÎUrth���uZ��}x�Ɋq�!xS��w��ƪ1�;~�\ʹz0!+\ʈ���8�S�V��X��.�P��]�+˗��#ړr�Z+RAا�S�b��Zm
<=���H:�=7�[�`#��K1�a�`R~\,߰q�P��_����%���� �н� �?��y��f[��rk3�nu/��M�7S�<�V
�x��~Gt���e����F���PX�@���klEub����Mx��	OȬ|\5S�Z�Ux��B�13�`پ$a�FЉ�W�'P�N�W+�Z�<�W˟^�+����Ч
z���J�����L���U�ܘQ�F���1���.9�ؖo�EIG��hd�����t�&�Qu�[�&W��e*����,�-\�DH��P����-�0������j|L��֠��+�_Y5������$7�4 �AD��lj��.~�\��v�6N������fEQ�����Y����u����c\w��'�5M�=�J�j�MZ�3���\�D:�E%���`�@T��v/S1Oqm��B1�:���M��T��߽U(����\��=D2�cOim_��A�0-�c���@�욋�u���(���l��n{B�%�/�����j&��x�B1t`�˭,�L�Aϝ�c!Wa�b\�Z_*�㞥�Na�6-N����Zg;$w&v����������Q���2�RK�*}C{\�@��̽�/��J��e���w�K_�$�X����o=� ��m$�g�w�����{��<���c@��)�ܴ����
��V�-��IOe~w��1o�v�$�˖�[y��[�{Q�8=gZ]���7��v�CGry�1�T����Uəͻ����E�L\(��4}Y��(�>kdk��jl� �J�U��Tk_��x[	�JE���`:Z|�\��J�����	E�4t�Y��E�eh���eл(k��۟䱑��C��n|B�����ݷ���)���*eof��@f��5�i� ����P��X	�Y������> 6Vݜ8sްCr�"� �ѕ�%'�`�Ԓ�x����K�0&�X��}�.i/z��a��C7@�:�	#��Oc%�s2�'$(�]�,z\��~/ʌ�6������5v��}C���r��7'�-����v8�U�[���X�����7b ݈>���)n�6�7�S��v{�c�O���`}��� �����S�ȏ���i��l�7l�(`Uu���)�T:�m�(2�F+	�d;_��ۢ�����V�kW�T8&��q�j��c�nRW���$�5l*m%I�ޗ;�۔���s7=������o�6��$����Ĭ��s�ԹF��ּ�	P��N�"������RtӤi)Ee��o����ьA�tb�@��*�����ʺNE�.�_u aDG?�3�O���n2/���e������2��s�&_�t�C��9��~P?R���'ڍҜ���O�%{����T��5�-M�'�j�4��j�:Gj��`�	���4)��%�����O���+Jn �.x�/F�+ K��XRo����|CD��!��vt���,��W5�����KR"O�nZ��/f\,�����^���SDgVu��z���Z�Ы�����Ę�\�ܿx��	x�T)�)Px����H�K��������
@n+m��[Vk!�p�D|�`�w�@[h���u	 /��?W��B���Ul��d�2�8w�R:H�
�7+��q:�K�� �gm�_�\����K�7e��-[�� e!�����tC���`{~Fǭ�Қ�%E�D#��-w@����[!v��`>�Ӭ�����yM=�W����M�   ��`���I�
�L�M���"�BJO�L_��5�1� ��ӵ��T'���[��#I*�7�:��Vce3�w3�m�m�[� �8?�A���E�x��[��İ\���:s�t_�5����5W!sO�O�o��q/�y�s>9^��=���d(n��M����p$��t�gS�a��3���ZT���8��^�t����U���|J��b^�2�q�*���*���̩G�rd�|[oI��w�Cn���g4 lm��o�{��&�R�P��~�þ�g�:��D��|�E%�ĺ��7Uf0��������g��ŜA��_h�U��e��W�?���z�p��}n��,�wQ�n��/qO�5��ُ�x��A��C!.�ҝ/VMЩs�;��H��ř�T0�jy�����/*�P~r�d X�j�
���b���V-�� +�[�A���m�iQ+�1��$q�g�_=;�KC���w��� 	{;�JjM'6&��q0TZP-��[N�?�5�_�^�e��������=����ei�O=�S��-�����ˇ_D��*�a��T����[{�kU��ٙ���Q4J�rZB_D��}��r���� UD=H���ѢaYD"r��10��|�q��c@I�F)1/�������d%����ɔI�Z�9/6�pبh����4�y���c] �sF揞ž�z���b������~0���0� 	�aL0!B�9��v���1�Ǳ<oG�� �=,/r+��=�Ա+1�q�^���ԃZQ�Գ��\�I�v�Q]��L�Q�\*�[tk��*�ىgt]�ްd��I���Q:~=�T���W�Eg�/E�����/W�Ի}���fq��SD��� 2%�(s���X�)�#����(K��K^�NpU5��ђ~�F����נ���2�v�g��ȍ�l��3^��ZT�2B�XQq���Je7����GIg!�SD�_���ڞ�4,��X<����j7�Ԭ?9�f�����{ Y
�>o�ן�G��!�[�=Hmx�%�%���<�����f�Mf�GA�?���೓���\#�7�ځ��С|�tن��Vt�"ө�=�T���S՛���дI���׼͓:���G���뉴�"�@%pRd�m<tm��{ڙ�&�y�t��٣o�K�9^TTb�4��/���(����i�O8�ߦ|%O�Ej�0E�����gY�3�a�/��� b�/
4�[���;�	��?���Uu����n��x5�G�J<J8E�� �x��핕�	��v���1͑�,f��
�3�E�e� ��G�ܝ)��Gz���=eL�0z	���S�|7���ݲ��������ǻg#@�ȝ���@�ߪP)��aШN�����W��+f���w��Ӫ�Q�����#?�~?)�C�ﻉ@�P��\��9Im���fnn��
vg�`3=��y�գ�����Ǧr�{M?�V�a�;�" �;2^�Pб�+H�������@:M� ���SQ9�)5k�o��s��_��� m���ߞԚ7�m�9T�"x�4D���C�V/K�!PgT�ei�7��I{�i��P���&�Dq`��t|�f_S�/A:�'��`��xq��q�^��+���鰲�"<{��K�rt��ڻ1d�-rm::�t�Nz�?w=8��c�맋�F��D�`�[9=4�OM��!��tR��/� �Z/ͼ�����4y��db���I�BS��M@0���'�ԟ�)2�Y�d�䏫3�'�a|$hT�/=����G���,>���+�%Q���͌�=G
�I�۴(��L�Mu%�n����V�=��<���(�Q�Eu�!`�?[�Ѵ��˻=r;uY�T��gO������8���G�m%[*j��'�%ot���M�6��Ĉ$���8��l�"���M��͉�.	���5���/L��Y�{�)G��9�	 (Q���.�_ɂ���A�@,{p���mP[�\��N�a��~<�}��N���>9�����XDYw�-/g��M��u���6���8�iv��d�ա��pš��
���|b��:d���C��K��I^H�m#֪����9U/ $<�^�i測8���4wh>bh����W�yj�]�3I.ߨ�+sn����O� 2�BTxW9%�*G���?2�	�<W+k����ِ�g����8�t��?��^�����Œ��é?s�8����9��b����RZT
�D$����ϵu�"r%H��P�r9�T���c�J:]���Ǽ��UVƜ�8<��������G���ˎ�{�}��� =�������O�<!��*[�ch�>7��Kx/�uƀ�)	�x&/�P<Dw�ef|�A�z�ȴ��)!G���5�s�2�w�\��"�<w��΄E:���D#�}·��ӡu�2�#����0)�#���p�9g,���KCB\t�SS�\���O,��f�����6b�X��c�;�9lĘD(�1l�,wv����b��v��eZ��^ B�'B|ק,�FĤ��ʨ�ʘ�2ܫ}�ع����3m��#�I�8���,Zh3g݆̈́f��#��2ͺ�t�i��e��I��)ф�
��h�+ �����������,?��|������u�:Km�͂�5P�����g�:��9���~����L-��}��{�{[�k/�S�v���,���m���|�	3^l�r������N���
����힞�@t�l�wT�GG�a�s&��eUL`�^s��oM��µ��b�� ���S��U���oo/R�]�7 7:�ǾJ ��~�!��K�����W֍�<l�jT5Ru\��4�Qw�>>��B��e�2��9��2!<3��<\��M��<V&��&���erhڠ��5�Q�H�ٺ���'M&I�1gGhT�|����g�;ɸ�D�pe�J\���u�"C�jm�A2�O�?ZZ�r��nm�wbڪB2�⣓AaJ���Y��z�&e���A��6�V�#��
���G���Y���L�[۬B�h�TiM�&���ov�٫/̡�*c��ڀ��7�����%���@��r ����k�s�&[P<��R�Ju5��[�.o���'�����N��u.jX_��ߔV$ۓ9�i=G�a5�u��N��0Cy����<��k���櫅���h�8򿯘^`�}'�������Q��wⰱ$�~A�g��C#-���q��?C���X��p����BP�+!O��&���?���sڹ9k7���y��$��pc��#�ñ+�G�;�<����F�>(�}�&t��������	��PGd��ߞ����ߟ4s����i��i��ֳ8��$D)ژ2�ӿ�>u1p~��V��{3ay�������*��������>���Z�o�cjY�����t����˂ǵ֏��y��?ҌSXҜ��@�B|�R����Ь���m8���ܭ�8[����ʿ�z����
�i�i��Xy��L�S%��@���. ���/�������|%?��{I؊>�+��ļ/��79����4)�o(�lN�O��ī))���H��>n�p��clZQ�Q%Iݙ��U�DyT�mE�LLt��iIG��N��De������?���/�x���f{i,��J+յ�?o�i3��:/-��U��s[پz..���[�dZ�(qQ��Ci�<�W��f"`+25�AEMO�r���|����)a���o�3���f�R��1�f�nɮV�d^�����ty� 3AC^j��9�r��w�d�����e�/�9`�O\ο�Җ��eO}�;��[#n���^j�*o��f��0_A/G��4z(���ܞ��I�L��O�󈔧8�&y�0Y�;��j���[x�Ș�./�U��]J8U,�V�8kz�AA��D�
�u��2u���L��~{��V	0! Y���ͪ��<�?�I )ߝtx!�����㥪�N'�lIҲR
+<
�p��3������a׫����������"��H��A�y����J@�pϑڹ�r���Y��֠��Q��\	�_��L�N^Ș[%ʘN���j�}q	��;-I>o�c�h�G=��(�}��^��^�9xV�⢻�^#ĩ*n�6�*�w����h���%�E"/ GO�*WB^��+ݶ��(� �%�y!���K�Eq��qmc�&�61b�>FEߍ���"B��|�u>�v�����S
(��H����H�m�j�Y�L�L�
���0O5��Y2�~�H�*���B9�����\��H���	���3)��uѓ|�U󠲼"ҥ٩�˼����h�r%'��愤�u��T�8:����g�������jI{��	�����a,�b�H�V�>�~�Cv�T��siM�i>Z;汴D�t�Z�S9���~IY�ѝu���D�*�B�����0ӊ�osu��������o�;�\eΌ�R��k����"�|>cK6	vn������2��y��9y�F�{�#2b=u�^���@6�����;�'����'ᐉS���zR�+��w�K��뼏�s�͡q!���tdꇀ�z=ݣ���k��:�ך��/�]��7����e��4���֏j7KFEf�u_��л����­4�*m������U�c)��5KdMX�^���śz��»0���@���ZޟY�/o�Sw�#iGq)�Ǩ��Z�D޶�g�@�7a�C+7vUѤ]��<I��^�������`��C�w�7��v���QV4�zFY���8�2<� ����:�鐚����k���1Y~������N���&��_��ړ��{!s��~k6�7ݐ���F��"4�ҏ:%���aá�`�V�c�R&҅�';�����������Q�m��Մ"ם��V�M��ևS�/�B �9�s�
�bf!I�� 5���U��;� )w�>�^�����tН���)r�hԣ&��	�G�(�c#����Fk���Z��� �9K�Ĳ((�n��LQ�*��.��	��d\?�\��U�(��!I����'�05�_7�)�ᣨo�4'�2��wn��\f���3���׭�/�� ����5{˭��`��a�Brq�k�'[A\֥iߡr���l1���H����UD�#�v��!�%�yJ�Zz�e�n8��h:�T��[����w]�R�M���Mv��Z��_�l���v��������O���֝k�yͺu�U�I���)�D�m�aL	0���wl�M�m�Y�%[�Ճ�+)���	��E��fx�5��n|��iR��j��t��D\Qv��Ez�	�3�U9��^���<e���t�I�A7&��sfXs�'�z����۾�:����a1q��ss���y���~	t#viM-�I)(:P�Фմw{���Q]>�vW]��:�[>/�������C�6CȪr�r.�0�׵���fM�n�d�ǐ� �3�ъ�c�a�yN�����`���fKf�WBx������JٔB[�E��if����(�Y�L�A����~�f��m�Tu����Wd;u��ܕ_?+�Y-��#���2д�\G��(O���uĤ���>����2,6ic�q��$�g<.�T� �tZ� 6P�۳���(*
��`�Z�m�p��UT�^��~��Ɠ�{�7EB$�%b'��IT��:���Q2c�t��Gx��@�s��8x�Nt��x�����p�����=�1>=��ޞ�/'ݻ쒒?G�����2FCfح�ҏo���4{b�(�����;�u\��<G�/�	Y�0��w��4vJ�m����o\����}89c��-d���}5�b��&rM56����^o]\$�Pҥ��s�I[6t]#Z��0��:�=,;��Y?�� (�VX�V6C��>c,jx	�����5��|v�/�TW�U����b+0�b8Z-��]_m�![&��_��Gm�<��T�E;/�x���r���N�9<�g�f���U��%o���������U��"xWI�D�q�w�u��ĺ��,���#Bm���NE����du4e��d�<�\~�02��\N~�`v��RA�=S�P���R ���X$|~�ѝ��dc���S?0�X�U�$�{[q@���!��~ɀ�V��R2O�1��� �?K��XFM�ݱ]����I3O��ff��F.�Bq�KG���J�TTH\̐�g�`$�U��S`�4T���]�m �-���D�P���v	��S�*(���n����B�f�=��Sݥ�x�̯�+�v�sw�&D��
0������,�������� 7��&#�#�S�T�۱���:���q\*�gp}�f+�|���>r���
A|������:u�!�w-��m!�O�ԵvKP���.&����P�D	9s��z'bzʝ�CN�-X�Ѷ8}��'����
�u�*�_��K�<��"g�#���]# '�2\�r=Y<qz��R��i�% �ơEױ�<#cUЅ�x�*���~�5"M�fN����z��j���h�$���M��H6&7Y��I��
W�؇��� ;*�c�|�4��:gy
�d����	�|[�)!v�3 �~2�\����˝8y����b�"��������-gug:�6z� w�Ա����?�rY��HQV���~Q��
f肇�Ȧ���a�ι��0S�s`�KYK��ZR�6�dS<�{OZ����f;j>/HZ����0�O�.kxE?]} �w�;�*��Aj
m�x*����"sܧ,+�:`Q��|�zx2vR(��@�_@%�kb;u˻@���ה�!���|�­K�N���o�8�a>�2��Go�:Y���E��	��L�U�lp
6I$G�h�sk/
��T��|bU�؋8ʓPn;[
a�TĆ�M��V�R�Tb^�ܹ��C`y����ӓFS���W�nN��K&L�J(~H4�m�Ú�5���rʤ��-���^t��IXlV?��I=b�h��M���X��A�;����}Yi�rm�܉���i�1�p�]-�k��iK��~@ar���uk����b������|�e�����|c�q�Z���R�O���fA�J����{K+(F�<Yǯ��5��"6��n"F��f|-͗F�v6��|��Ǹ��/EzU T��ts��O$X�T�A ���Mi�vh�Y�F����XN�6��a��M��7$�)KM|���)��>�M����%!�#���E�+�\��$� rb*���D�ߊ^d:ս׈Lz�'���{ yѶ8i��>�H��.�,	6vV�����w�`"�Ì��k�����8]�F���ͮy���7�ެ�L�v	B���B��ebq댧e�N���J�f���wԣ�b�����7�m�;�n�|a�y��R�;�#:V�f�;j�s�������GM��I���K�gޏ�^��4e��I��Y��B?j��"2�;���!F����{�.>t�;תRT8�T8�r'�B@�[ZX(O����B�g���7��u�QhP���~�h��XsN{��I�� ��KxE�@o�|L�9���tiG_�F �tp�<���[$�:��6�q�ֿ�k Z/{����� h�冄h{cf��eYr)�8إ	f��B�;����x��A���������T=�&�V�f}�$�7���#��;N��ӎ&@�3o��$h���̴>i��j�B�dJ��8죻H�f`.�KP(��<����g�_�U��"��Q���o$��\��Fk����s�h���1�ͭ��o���T����<M�/���C7�&�e�m�?-�o��)�����N������`ͷ_��G{�ȟ���.ɤ�r���CZa�@����{�o$)J*�%��j��~>�[���X��iO�tr�~���o�R���Gx��\�.R��
t�,�C;��v�ѯ7�6��2[љi�	0�ނ�ȐעQ=3D��	�bۖ�~_<��Zqg��R�C����=;��PQ!�h뺩�|��d>3��UP�z��T<�rI���0wCxUC[�S��<�dKo��]��"���fm���%���'V��>Nr�5+�����_Uڗ�zaL��D��-�$���$J�x�/F��,6*Z�?��\~P��2�����LZp�ֱ�'�<_RL���00�7����Y2��!��B���5ǽ%���5
�' � �f�g��1A��c��E���l$�-�mך�VLT��������=�j�<i�9_�3s1� ��a��u�����8�$�-��t4�N�o�BG�$�d�{���T+����\�Ux{�k� ���?�a�p2���s}����ʍK�`��X�Q�����w���ʧ�$����Q��+���b)��a>�P����L��ݫ��W���%	
��(^Fg���o�VÙ[�^?�|gWjK'�) 4}ۦ�<��M7��+5P�Ξ�ld��qm���.t��\�t���cؒ��݄�Z�z���q��ѯqב��]���L�BKx�w	t����*^X�c;[�r�R]���V�̥���O���_ql!�s)6��+��Z�W�Ȼe���C>�uq�W�nso��@��4�I$K	��xZ��8h�b����8
����[��.��m�4����~ש�^�v��y�Dv���i�Ӌ���_ �`L+�H� ����
�TH��;�Q�%`
3>���b�Lz�y�B��|t�8����9���ד�O4����O[{-��"�+^쉭*U�.�R�3%���.�J�?�|�$J�a�s�M����f�cI�� M�w������_�n }��`��7��-5���Se d/�����Z���~�Xjc/��gb5�m��X�
�W+P+*l����*��çF��'>	�`-�I),ɴ��9*6�P��ԥ;"��unv���	��,Y-/��f�M�8�MoI�?h�Ț�j^1�G��.�6o5���~e���'���i���ĥ��7V�;7]��Ф�<2�f�G���;��C.e�ۄK�v�$i��������{O��	2;�s>�?� ���Q!@�5 zpq�K=��ÿ?)z|��W�-T.�ѡ2�ZS=]�b��UpPo���*̐�9Z-Km
�(��{�@߶;�]��9��H�Tv6���)Y����O(��6���p݉+�G����:�߻��7i��h&{щ�D��{XӦԐ�䛓��+�����Zam�lSV�@�����γ�bDB�>�a�7lڬW"�Kg���:���R�vL�����.&R�뢝i��H`)���绍���}�?�s�W�J)�/�lxZi���?Q�*򏢯W���,r�2n~/��]]�����kJ[R�=jA�ѵ)�9��v�L���3���
2�Ih�kƠp
��j޼����p住�4�zl����&=-6�Lϡ�����N�}�q.�E��yM��0�%��&�,�x��4n_=͙����c�-�3Q")��:;���\���JU����q]��m�HOSSQ�����e\���@H� ��Z�M�/a���n2���k�n|���)��A$��ag�X���g�{՝�,�ƪ��?x������H2���A �[�cU[Z��գ_�����F�ă#b���R�	����r�Ҿ�|�Z��;/iZ��e���e4�*���'bЀPb�2����U�����F[Uh�6\֯�>��V�>��Նٛ�h^��X�L`�,z��3$�R�,�ŝ�Hk_�e�B�8p� D�T�����X���� MMf�v�\ECٳ�S����.F�.���@���D2ӱ�e�^��_��ӳ'P��E��t�e?�9�rU��ڨ��a!�����*��-a�3/�}���c�����`,*D"��Vi�q���R�G����� A�썶�����M����jщ9�]Ɍ/��^V�1����zj��-�Z�����[J��ǺAZ�,�����ၦ�)v��,4���Z�̫9�&���[��LHs��N�Vǅ3��T��Rn�����	����",�3�ׂ�|���!!�gS �ُ�i�0������1���:�d�8�ֵ�d]���t,9��=�tU�� ���~3�0��0�'�����g~-�rS��F2L�Rۅ����cP�ί50��j�b�c��C��}`#)��-�~��n؅BpNA�XI�7��c���[ )�X
���U��y�����H��Ӥ���Kѷ	Z�
8�;�^��gZ긣�8_�����V�6pq��' ������u�]0���������k��R6۟�K���гmD*�51�si�R�s�J��z,% �#�|�喹�'�R&A0~Sz��������M��l`�i��-�g�ȶ~���;!_@����*����=k	�T
�n��Sa��XҤ�9����k8w�rR������U�$W��m+�����1��G&�喆����� �Տ��'�j��fKc�CD#�j��
ba��HG�UԔgҪ��Y^U61�=3�[\,��4!1�]�H'ٻB��DZ�Q��]I��R���6�`�OHH�U�;�`/^{��̚�w&�g�|H��<�=:PA�,�H���f�JY���12 ��%�����Ӓ#������HӳeݎX�3�k��u+f�x����������"�Y�v/+Uv�|XH�9}X���y��M�$by=��Z(��*�%g����	3���{ :��~���L�΢YЍ��-�2G�S���6�]�� �G�����<��
�/k�o5�u�v~b��MU�9%;=s�
M܊����E@���z��D�\b���;��[��#N�l�L��/�����[ !��U��!K���y�+�V�k�<��׾�=]��zs��V��?��^s�^`�P�Y�T4�'��b����]|TW�.����Nw(*��'���)+��젥��IS�p�l[��Z��E�jy�|�db�d~#��f��g4"������x^�Z�n�4ی���s�kV����8��?�jAI։��$z-][�䋇�g1|�^Q�z�6���@�����|f�S��|�?@7}_�����~y����l^�ǃ�G�~b�=�!��+��m������&~/{����<��;��G ɥ��b��M���N�S�^��1��X��/��˚��&�'(z	z����m���׫�}���UR�QZ��>��<�'�c�"g��`�黯Ǯ\)�sJn�oB�e��-!k�s��I�Ζa>�R6$r}Ssc�Q�eU��?ڼN~���m�S���2�o/����=rZ�r����~ �a�ލ��-�-Q5_�TJ���c�Ȯ�Z������Z��l�S���x��L���D��Մ���\�O���]؟�|zw,>A�T�6=�.gc����f(	] �����Hv� ��ޤ��J��E��fK�6y�&|�4�q=s�������� Y�m߆*4�2˨�WMS�p�N��/@�h��恴L��e��̿OD�h]\��C�6�|���1Z<��ֽ��mӇ�1�1\l ~�n<���/���~��	*N!�W�v�7����)Z�'݆e���v�e�L#Q�)ߎR�Bj�K��}<`Ӽ'ô�F�4tWTm��m!��o�BK�\Լ�.G4�̂SZ�Ul�2룁"�nR�#��'o�i����e��&D~m�d��uW��K�h�kip.�&Ɋ-D��]EIy��H\hg��b:'Lx�l[uC��<3r�}�y�V[x
�l�~��l�=w���4[ev���ث����UC��R��5�@E+w�@�?$]E�L@��\\%������� 4˦rvq�3��
2Q������Ֆ�8t��!���My� ���8_��`rISC�b���J�mY�+��*j�����Ҿ q�p��a�x�~w�1�yQ�?	�92n��@�M͓#�u�"�����R9�Bw�$�M��_�u��OEҠgg������J0^�4��� �>w�P?w�`:#6?[^��a���՞���k��z0� U��q�1���
����[�Nv>���3RRJ�g������|'�|�R�!�6i׳l���t���.�p%L�/�_�V4W��^��R�ߋ޻~�7eP~��(�9�x�m��;?_O���?��fwl!P���9n�hu�Y�oښ�zC��&�r_�aɵ�3�T����ZD�6=0�(2{�~��XE[:)��6a,���t������Ĳ��R:�U���Wy�۲}�y&>h?n��'�����������>�G�<�����N7�f%!ݓ|N����۪{�#8П(w|��2�4�ivl����;5�����\��u���&�݂�YR��j���>�@'L=�������q{�j	�y��� yz��1�I�we&)^�E��C��a�?��`Z���¢U�6�������gۊviƣ>��Ρ^R����Q���ۀ5�%��n���꡵Ӯ�l�/����%<���!/)��s�:�p���)˚B%A�͚/��wN+,bip�ݻ�tm(f�ͦ���<��e���<w� �:��V��e۹�o�Sщ: :=��Bn�9�8K��C���}������zU|�{Q��4�v[�?����v�f�� nm���VlJ�>�xf�g���8��m'���>@�>������I��D�?o�-M�E"0����f���]Ђ���|�wAX�ϣG����^E����&�vN��3B�ܼ�k��~����y��˄ss�%�/!|�v�@
���8
�m��0v�2.į*�� +�K��F�[�mcj*W5t�%ZO�P[ X�T����Z��d�v���<��. �����"*WWQ-i���8߱+���-�ɚ��Q.��pyh�Mwh�)�UP*�Λ����e��H�fxxF}P���C�nO�v:�-Qv]���1KQ�+Sm2Q�m�������&x�O�0��|�i�͚�pD��8�r����_����5=&��	;g�m,�O.�q��DŔ�C<+�.7�7y���z�fr�qM��Ho�17ߢ9x�i�q�+�:�0���U�L���nM`�P\����mR|k(���&8�ڐ,L����o��}\�}�ߙ��|����v��Yd��9E5�xF��*��^��깳�r�[������ԍ?�;�B�=��:��u��̜V	�k:�Dg�衊�3��BӲ���(�L��n	���~���+�����?ۙuv�3.���=����M	Cо5\��:/8� ����}A;��ӕK6���Wy_+?ESK��IXY������e�>�۲ܛО�k�_�[�Z����ö��Q����,�������}}`��Ӟf���ᡓ�fr'ҡE�	Y�\��֑�i�P��)@	]��L��>[y��휻{Q�7	���W�g�Υ�^AK�~�G��%v � $�-����h��m����P�b��M�N���`9pK9jL�,g�w�{�D��A�`Ezb��2�|aA�jw�*~�v��E��ֆe�)<����B\5�����a
b�nbx>� 4�wH	�ϊ�PZg�����r�|$��
b��H������t���i���z"膂����?������O��R�|��٘��v�� �Z�MUI��&Ԥ��+����{g���3?:=��H�OB�9	�Ƌ7n���[�Ԁ�BVa����������T�0����pڬt�/�sy�ה9`_���I�zK�w���5������*�4 �I�B�xS��:����0�u�J���?�m*�a�Y���&ȧ�����tUz~4LIp���7�����k}U|��Q�����߁�'��W�U��=��UB��o�$^�q��>�܏��c�-XK���`]�N��B�T�ϙ�״nҢ�夳��`՘��7�h4u�2_L����ki�S�>@^����\J���δ|F�����ʋ.'3Ր�	**Z�
�m����vM�����vLdM��7��dF骲ń�R_��G� �G:�@E� �O� �l�����]��I����� �Y�	��P(�=%̐1�|N�2�L프�'��^l�c�8ːw�X������!��:�ͣΎ3�N�G�����X�ѧo��-K�7��a��y�� 䶔��6_��/�h.c5�êh%%�|}ȁ��|���������	�(�_L���F)�������|�#.�G�=���C֙��r{u��E��?�X�o��%l��L^ە�m�ܐ��.����X����?L|TU��EZ@�[���.�i�n��[����t�tww�;W���YK*�;{曙��g^z��[�Qee��./ء�������[��б@?�7��ܮ\�-z���-�s�ښx�/:�/�f�&�3?�"���U�|����9q_�L�z7ű�m�W���Y���Y����#����R�ѷ2kH��ܽ�_8k7�ռ�ʔ|�P����*�q�)��}4Ë�Ɏ��c
�՟ޭ��J���lwō��sOS\�V���9��XT�y��%��)�u�,�^Z�Ը�s�ѥ{D�D�z���<�f%���́���Pߟx��S��{T���z/�[/Lu5fo^u�k�c�G�^Z���o9/�T.i�m������"G�:�5}ůK�fF�Dɥ&���۱f�8�f��/������h�z��W\�H���I���	��P��g�*E?��
��j�X`�rXY�m�t/�XQ����'��cǸ�i�
��ԏT�'a2���)j��1u�Ύ�$h ���U�贵�ƻ���7
�Υ�^$F6'��I�Y��te�W�����@�$���u����^f�>*N���eOn���D߉�����֎/����6��3 ;\�ҧE�k((�ʆ�3�
���D�l�e�s9����3+l ]��p���� ��^ဦ�D)���]�lZ�w~�����yx��V�t�bB�棽�����%�u!^�TO<V_/$����
��M��υ��]�(��z�S�~�|��`�{�C����4[)�]�7�H?$���Y�q>��}�x/�p7���ְ��4���;��Dk4��	
L�T�n-��W;���j*NT�xd7��Z#����k�#	[!�7��L{�~��u�L���q�_��j����I���A%�ުc���\�η���A�4������'˚4$�I��4���R	���C J��l�4���0�ܰ/�90�N|{U���ü@�����ު렞����d���+l���$��Zd��S�;�����!��qM>�wa��c�и�)ԪG��6�u��@r��!���
v�ϑy�K�.|����˓�=dn�Z�U6�i��zy�,p$;+J���#i�WK�<\%)48ǳئ:OU�-� �斱r��sʌ�]i�$�K?\�:YyC*GчEK!��x��ׂ��/���Vs��R���ނV/9�'&t�8�D�喼�H��,��s�V���p�Mb�&�D&3��^r2x���:�*#�{��<�z������>�oR�8��ϕ�TQ��|I,�j��E#�Ҙ���>��I����ބ	s�Q�Fyw�T�H���������b�QҾ��i�ceC5��!P�T����\��;Ώ�b4� ]��o��&ܚ~N��ՈUѯ\�n�N�D��ߓ��8�����Ќb.��^ ��o逰�d�#�_����!?%�q���+�ګ���l^.�6�^+1���>��)�b���ؖ	�5�E�1N��~�y�`��b�:�@�f[4ԓ���T����9�Nh�.�a��J.�'Os.g�����ŧН���@�T�����4Xx�X�x�� ����J�Z��7�%�a�7I���	� \��S9g���A��H�����B��ê�d�|:dbb�'Y��Uy1s(c何Ղ�$}���1b:�Y����J��%#��o.;��a@8�#
QD+�|����ӳm�&�T�"���	�NJ��~�G+xq�|:���sD���&aro y��r�/:ƃ���]:꫶�$��"���V�����)M���jl��E^֕d[eRց@{� �_�o�����q*a���M�&.6�h�X� ������	|n7�!��u2��K�1�Um�Y~�+���t��d��v,��o��0L\Sr��s��|yr�}��$���7���.�x�k,I�a'�k�9z�D}tQ\ej�K_X���� ��c���8���1}'���7+��z�.��`ʨ�F�pl
�?�8]u_��t�(���.b�4/?cd��|���դ���:e{F��0oo�Զ���	Y^�ߏ�*[�{:.;�v��(��'�a ���ŐN���7mE԰|����ކ7��~�U��S�m:��\".0��|]NH�s�wY�YL���i���"���	�a�&/i�,�@^q��)a��
�=3u�����.�2��H��J�A¸�tFi������ �i��u.(B?<��o�xp4�N�0 ��0���I[^��
�0��rʺ�/w�ç��/*�,q��wL��t��W�AN]���QX�VP��E}��������D8�G� �T�� L<�{��W�����@˫�ߠ�s���{�l���{/7� �xt�GD1���K��W�{v�C��3rs�(�/��vxM�rC0s�Jf	�Cd�kJ�@n�.2(��R��PMVצt
x?$�l��O���,d'�_�	Gܔ$��S�8�畜��z�x䏜,�vy���?y�Oo?8Dy]*YlM��,�E��w�WwRJU
;)���+�}�S�h5t�b�IGG�%s�n �!�����z����%�����$�sI�� ���������kh���Yr�B�z��"�=��xL�r�@>hJ|�[�4���Y�=��2�q\�M	Sb�Wa�ZJ��?Uv��vJ.�]3'w
�s�<��nVM��Z�=ǿ��2"������/���Ľ�A��e���n�4�eɥ{]��Fo���=�3�ԣ�VK� L��+���*)���5�b�J`�^z����_1�\LN��EY���g�AG�"g�輽��rUG�&�:������,��FF���0�%'vM*Z����4�D�:�Y�]m<����bV��j@:���Ӌ�g<^��3}�^��l
�s�A��R����LNA.����ޔ}���Qf��&o�m����Jhv�I���$��ʢ�B���![P<��4����ᅪ��7A�c4�Q��O��.�5���� 2-�Yى [�g(YVN�Z�t{ܹ���A���,�xc<5�
�}�"@Ѐ��}׼����N����86W��N\k��}���T���V�'A�}�d�N��[R�����x�MEM+�#�O�n���O���y	}�]��qͅ�o�g(�9
	ԗ������"�t�Yv��2*��i�@��V��zp-y?np��O|ͧ@��b���F����Z����z��������LEѬ�M��j�MDΘ���i�*>������9*�3��b���"[�\��sNT�+( DǂxWљ��ۧ�*�_d!E9gp�pOo79 7�1�~ke�����SU/?�X��	u�M���
������f�Dpb��E�&5�� O���Dܼ{��ګ߽Ƹ2��#�U$���ZPN�M��\u��������)��LV�c��<�/�\gϴ!J���4�f����!�Ae���q\D�+ �g��&~�
I>��Ⱥl\d1��e/Y@5H_�@���!Q�Yn/*�r!s�f��#P��ar�'�L�(^q��é�.d\��@�]e&z.L���������,s7���ʅ���x��朰��"�������}$��-��%�7���y�?�G9�D@n��5#P���BK����:�w�Ҩ��=�y�g���Z4qޜ+eY�e�,�M��Ю`��rnH¯*w!�1��=q�?��U��銧�g���]�b4�nn#}y� �ڥK� ���J��58uB ��l��a�r �_��r��:a��yt��4hB�����m�M�����.�^��r@b�&r?C����L<Yz�Cf�1@>��)o�h)���M�g1
|g�W�o����s�S	E����o`��D�'�
s&��q�\����r*
�3-��[��/ft�ז� �EtX!�W+��JlD���w��,qT�#?S��_�2)�Nv��\��a�j4�ݢ��*���l);��Q�[-�BJ�~�� j�� 2�Dħ��DvH�@}�C�C%��⮋D�q�Mg��Qɺf�������+�l?!���0��R�l\�0��a�	B��T����yŖCS�!��}��V<�O쥿{�r=o���f>Im[�ޑ_48.j��U�=LW�J�щ�7�]x@B/���chy��h�|6�;��se�U]ˑ��V�^me�/m�Ԁ�>��!�LO9P[5��6���x�>�Q��H����}�� �}z�� �9�@㔥��^�1z|'�-��d�"�t9|�w�����UD�Y���+,=V�ͩaQU�~�e�U��>\yhZ7�<��p�0w�Y��I�����l���s���j�dp�j +���\���s���J:6��� ��mS��<�N7}$����bC�D�]�������-y�x��Y�C�GU���Uҟ�Z��x�]ŷj8��A}���C���o����1����/\�t�*�_ �:���hv��F�v��*-_�=��? m��������'��%.}�9Sx����;yQj���%���>+���:���3�("J�Ɲ<�ϻMi(���`��Y�Q)M�\�[�&O���z��[^�ڧ,�\=;�^L���2��P����V�Z��Xǒ1i��j&��[��.x>�!���QmŎ��^=O�<w_�˓�B��>[�Bn�~Sһܔ]0:<�:�R�(?+�0��UVJv�l��j�b<������
����}I���O���ڃ��O�[3��q��b��e�SYZK�����t4sv�K��`�b�e�ʁ_��Q�+�m��U����f�P�2˽ߓ����bLm�&��EB�>j�����jv����!�F��\:��3<?;�E�L{�1�e�p�(�Z��7��%W22���WĜ_���jp���p/i�̻P��j��}��I��u����p�"�i����iX��:v�pWrS�'��&8���6Bf`��+8��u�쥽"��)�$^�=�N�g�N�2˼�b>�QM�Gװ�ߊ�`��)�|�!9��Q�1�:�Ι�[��~r�7�����tX�9/>�9�Ic��9R�T;���^�+�-u��Tal}�]��ݛU�7>����]�~ۧ��˃[�@7����ݍ.�g=Dq�鈆�u�Q+z���am3�QMo�2� NgM��B0�&����e���o^�fN�q	�.ٿ`Ŝ�,ψ�D	<���ʒ��O�!(v3�y��̼6G���k9a�.��y�q�d����2�cH���	����O�ˌ�������ٹ��D��ч�'�y�ʴT0�T�'Z�\,�a?m��t�*ܤ��g3Ok�Nr߹�4�M�����q{^��!�-�4KU+��0�q~���zN��tEˏ�N����:�t��&�hX��b�Poʈ
P�K�)^یE}䂓C���"?T�U����O�X*�f.��C�T�+-R,	�qlbR��hk�Vni��T�!�|�	�zVUH/.��
-�I�{{v`BuG�ح���9���0T�U��e:�0��/���IK�J�R۔�U6���(��WXm�noݎ�ӳTstsl,����G���:�rSE����D;�������H�u�t����N�z�l��.K��4�gD������I��ʽZ�fIJEd��E_6�'�1+}�'1�_�Ǆ+PHp�;�'L*&i�-�=結���?���&��n�z~k�bm�8Wr��Z*��Oܐ�%eNmV��?�"sS٫_��o|U_IK�����Z���� 塱��[��[�S��Eެ��#+M&�H��ѷw��g�l�JRU�T����Hd��#9~�:r�4 �5����f�(�ȮJ�����gl:@[��]� �(�9C�uKE�v�u�^pAW#Z>����PPl9?�i�

���R C_x)�O��oE���p�?�Y�mo6Ixzݍ%��?Y���q߸���c)c?ȯo��Z��0j��ex^�:8����6�!iE���ẙO����Խ�������
e�p@ҟe(ﾤ�h�7����,�;�Px��""��#BѲ�Tz�ca�DO5��RiW�ĩ^N�|�S�5����7����S�\)dz�B�/��1�ʵڑT��KI�лk�����p�,��I|� I;@��d1_X�����+���Y�;�B���AUqW�
'��&\8������?.��D�?=�A3Fv�8`&>~��4?Ì�ʫ�˚`J~J�kOo!NJF����%�����T�u+�w���\TM��c�kLs�@!O3\X$N��1� ����"�}����/p5tA�v].*���Y�h�jIk�~��( �����$���o&U��S(�[�,��1E�dPi�
疡�,t[��� ��.���;�ĸ�cS��""let��*s�1�ah_k�F3�h�vK��(��EI����N4E�U\g��{mD�:9,t=��b��N uZ���+)�M�^�L��mʁ"{]��Rֹl�����Fd/��3����=SS۫l��yE�,�w�Q�A��h�%�8�1>����^�N"��"(�^���%,N�����V;![MkDQ>I�~���,���M���oI��(�LRD�p��`_5�c�"X�����k	R��`�8�H7ۧ���+1\������3��������+fE^�ް�OI��P'�F:�0��	�� ,��}}�/(0)F��g���?���ۃ�}�5�,�Կ�����:�lz���s��7𢝽��Ɔ��|��Ť���Gh�����pUz���O��#G D�'\���9�H�b��5!��9�7��V}cxPw3�x�;�ݐ���ձ0~��"�� Y�$;,��>�N�qc0�O#�sIJ��N�c�71M�qVv*e���;�Y5��֧�0���Uμ9��*�]�<u����>I~�E�3�hB����.��G*�������%���ܡ ��}&QE�|;b&K�Q������Y���������}�:���GnmH0�u�e�[ͦ��b�� =`-�z���v��=����E�?bL��C@������$�L�˃o�����`sO���k��=Y�f:� ��L���'�?����c�bţ��2��C���$/�� �ۦ���b'%_8�(�.g���J��Y[�G)2R9:j�%f�H+#`��[+6C;,��1Gޡ�9���9��g:_�@1T�P�5�2ևJ�Uu1mY�]	�U�0�V科o��m�Au��(� xy�0������W�;T� m-������%O��ձb���d�V�2���g����v]'l1K��ʬ,"���n1	p��?}���l%�872�œ�ӵ6��_�����8�ń��BfݹNddRvĩ��to�����N=8 D��|�ݍ�
�0��L�T&UI�V��Oۚ���(b�"k�����//�LX��/fA�L��^�$��]�%�_Z�>I�C�e:ۦi%��@ESD��tL�S@ڇ��E:v%�k#��b5.}�o�j��_3�
��_c�9G5����F/�!�����p���>x��u:����#�2Q���D-K!�Ӕ�J@���R��]d�y=Z��$-Jy����N�"���ڨɴ��re��j�܊��H���Ȥ��?	�����AP%��i%^��ع}�n���Y�����Բ�H���g�k�5 ��3o?I�0�]!P�W�} �@����R;9�i<�*>�v9imYC.�3�����2^h�n�0��C������v\���`<��,#uu%�S�� U��Vf��#πo|5abW�_V]�'3N[�ݫ���
����]b����_��OǤ�ڑ���ox����G֍"v�+8?_�N֗�x���K�_���:������I����*<�XP��E{�RV��ڝd�0#��`z��vK���S�L����;L U4��m��n =�0Иs"~P��<@IU˕=���:����	�隠S٪BR�����;��}6��Կˏ�p�����8�/�������`�3/o��/"����G��̽˲����e̕�v�W��*>Uџ��2��|}�K�g��z�4O��^�k�'��>P��7f�W�����r-�ɞ��[ =�� 'i�ǈ�$�#I�>Z�kG�L`���T��M�1�W�$����1���H��������A�����*k_�����O�0��g_9Ս�bK�XgT�|K�܈sg|"�i��2��/{o"��.[�#��C�+�a�X���R�&0_��Z�Oe�fH1�'�i}����'Y���2���[��>{:$jF�T�M�\����6�~;�4�߸IY����D)w<!�ш��i@�@q��)�v���qi�W��	�74@C�'�LZԪ��C��<�xG�c��*Dl�s~�:H���<���P�P���B#��mA���`�b$�f��т��h5���f�L(��8֫A&$&Vn���&�'�1^�t'�¸��x]�開��krRI���}�~�o�5� j!�i�w��[��N[9�*8ym2���R�뀨,��sɸ�6YBh�;�C�1�\S�+{HO}�l
�s��C
�<I>�� ��+��=�zxw[�nIW��4%��%�q�u&���?�1>1��,�����j�J�k����\H��V�1����Y
,燌&"@����r��o �~PV��#
��2�D
�Mӝ�����A�X"f1�#暱�k<N-�~mҮa��Tz�i;=�V�_��D�ܭ��LW�4~)�"K��
�"."�=�������:f���Zs�����W��D~���~���v�:E9(h���즬�+�-(�*s	q݀7�XeP��Sw����,(��_�63���Iq�Y��#��}���~nJ�x�R����Ry�}�G�$�T	T?L��ZG��ן�+��5���N�+%��4�M�F��J��y�RU�
~i��Gڭ|�~к�n|p�i��XĽy�G��l;�Y��ޔ�}U�xxd��֦tsU��	����y��5\5�� ����@���t����W�@ �yE��j����G������u�ܟ�x��e�=�^]�?��c����J,W��M' 2.�����B�/��v�'�k!�P����8���$E�
��9G�ޡ�xl{Fh���^�l��ж��L5�9g���5�h���������@���^�/�F��o����X��O�U-'�tO2�֔��M�M-{�ۧ������H9S}t0C�AD[�|������&6�\���ᴳ�i���l�#��o]	���2�r����\nr�z�iBՙy�w|��W�?M��$$��e]��d�u�:�¼��$��ј�AQL�g��9�g+����/���fQ�]�^p:���Ӥ�a�q�zE�'tX�ı)�
���1 �a]�N[�ٱ��^��*�]<��Lz���38���t����T��%�vE��|�0(C���i���9"B�\��߭�>EΞD���Ee�~J�О��~ �a�<U-ϸ&����!L�����F����7eDîӍN���!ۏx�l�s�d1���Qգ��G��q.P�O�6��w��0B�m�kt��%�����~RC�	u�r���m���|�Ў��	��J��>^F�B->���5J���&^�B��b��6�^����ٖ�E��E���&�����@�h����w$B/x�q�G��k$Ï�H-V�9dkQ*>�3�<w���	 ɗ�a&���#W��	�[$��� =1&:��lh��	�é��eoi�v.B���J@�sjԃs�i�g�kj���<��Sbg��e�l�z�����`Q=�	]!��̗)aj�뭀��'���s�29��	?Ӄ��ԾO�lQҫf��n�(T�d.�tE�6�_�Iͮ,��kJ� U����6��A�p"'�l��
w�G�3�c�x�8�>���xtڂ�=ÒM8#K�|V�2*��%?
��粵�D�L:mDSf$��FF�Pֽ$t*`����˅;���)�s�	�N���ƈ�Z�ӓ��fWT�[9c�":r�ϳ�(]�͘�V�����磚���,�Ϭ���c�sg_Wj���ot,FM!�MB�)���a�Ok���j�F��{�ֲvn]���Uq�wWe^����B�ԧ��+UƮ������H�m�GB�X�qzSrܦ/���YQ���������jg�E�q�S0���*��|���l�
�+kIW8�8�u����(��Q��OH�pY��ߓ��v_��@�MD��f��G>��k�V8�Ɏ�n-�h��Tmkإ�x݁�xBnla��A>`9;]���F2�uq��㓒��x�~����&��/Iv"�o�I�jy�o4mg�n��V�e��ҁ�ד��/�����y��%u^(������u���볇�H�� �tłUM髞���+E������A��h�M��f�PI߬ڢ�����[�[=�W+��ʗ2�����k��܆+(-�V<.>��;�ԜM;���T2z�̬�7#"v|�k6>

�b8��H؃4�gr���&���kϘ�}���Vw�Xe���E)8��z?M�����[)|;w���?�<@g���Vr�m� �kR�e��f�=�ٱ��p��
)�v���[���]��}�Gh�H����Vo��t�,�r6�Q�fȣ�.�K��n��0/��`�U��pD��徽B�TVV��K�0�	0���J9%AΩ�h6)j����W��F��,4jC�+�M-��\ۨ޶z"Q��@F�ȺT���~��hK���9�㝥a/�S��}m� �-C����D�1s�	�)٥S�{�l�k$�C :���5�ڝ����'��
�9����Q""kr ҺTE{�J����̮�u8�jt(��;Ƈ�EY
л���\)Zq�',,����|����Q�5y"�op�5k�꒧�ȹ��<٠䐲��i`f��I�hS���}����A�c��Lǩ ����֩K�Nl��\�*��m���V��L=LV�=|ٷ���@[Nm�pM�2Q�w�bW՚�<!j��<� ��-�KNw�pl�����b�`�)���NO��q�U_�>(����d̀!ޚ{�rʥq@jZiG}x����������dK� �k��g�Y.��2�cGb�����]v�;��_#}���.�>;��c,�S4���vG=i��S�n����f��a=������<�t��rN�FWʄ��W���}���W�o�h�أ ����(�{�h=�:�h�����ϙ0mX��}��u^��BDī,	:�GG�5U�|sx�M1��9�������Y�|Ο����D�,vD �GT� �)��P��W���7:��ƑY�S��l��tV����q>T����t�M7́��t�9sK��o_�+*kqT?�9�~�j媮ʂ��y�pA�Ê�J��kE)ȱ[�h�,uD���ba�<?�$��g������T̛�)]T���?�gإ!�:"\�,���0�J��9��'���>�>k�k�?±p��{i���:�b��������Y�����l?<��3�2=�� ��׀t��ѥ@ ��ѥ���a|;ϥ��e��2��2;��{���k����ki2���@���yqV�4W&�Dk�վF��(b�Y�~(�|�Ry%H�ޥ�;�~����2� 2��yf��J�I�N2�h��A��=���TI~P	����-�T��t�>̊��4�Rc��g�4�[�[����0�@�����)�f��}*7h�uWa��.ꊏ�6`|7nR	��i����t:>!�Oh��Y�lx�uQiB�׊�;�C�n![w��jc~���I�M �h�b�u���|�S��8�L��z��Tdv�|�W�y�vMV��Z�)!�*���V�J����e.>ͽ�8Iz�^��g�/!Å$���o8��Y�BB� ~��e��_�o��3Ť��l:�V�圻��턑S[�X���_G������h���uAI�qmok&��H�\�$���T��%|_��̌��x�G���+Z&]�׋�������y�9m{���bܛ2>K6��ʧ!]�y@a���*��4��D_�N��E�) =z��,OQJ�� �}j��(e0��N��u6)�M9�����y��[�8�/8�掲�_��* �[����]��F����OY�
�u2��I��
<��,�&]�P6� ;��'���F����ˎP:Q�L|���`,�V]�0s[�DW�5X�d�r�,���y��.��W?¿���=\�H��5��=��F,'�"�%�C���J%.���
�K�⫈0F�Q�TKK���t5ty�Շ��<6���e݂�`���h �q	�+��o���G�^򜂍�=ݞ{���H˜�ȔĤ���������:�~:Ynh6�k+{D��ւW�[�B`�^L^ѓ.
Pz:���g�{��F=�#�§T�"gU�ٮ��v��@hI_�+�YqԳ��g���W�%�Ծɻ��r�e#�Q'5v)5cqj~���F2�o1(#Ta@P�ѧ;��⯯�E5T�P���8,���������-Z�8jn�6��y��su\�OK���E��ZYnϼ|���)�_Cs�& ��Zل��������u>DW��1JeT�)x�|�߆���x m4��:�Ae���nyO��0��� %Z�U�;�ͺmُ�f|��?�����[�?�p&|��P�V=8'�:Z�6��z�_� ��Z�D��s����������'B>� V|�Ӟ�b3�.��װˏ�LfW13!�px�M��EǱ?N�
1�������{Ҫ����>� S�q~Zd-"3h]�9���ƈ��J�-��\m�`�)�M�B�5��S1F�Y���NI���+�w�>t�����>|v���?RS���N�|9���6�����~Ǽuғd�y�[��c{{6�O�7�On�n2^x�f��6�T�V��y�A���(��礙���D��]���0���f�J������r��UI����E@x��dn4�&�`9�K�$M�-��O�Ow�eg;p�Z��� `���7\��hx���U���px`�z�!
��Z��4͠YW��Q�P���`�5/.�}�������q��i�§'y�s�(�� �)��F[�\��ē�g������-�=Y�7z�+-V����flU�����\|��{3-.��w.�u���B��i��C&�V&�����%��͗���G/|��+R/��#[آg1ޙ//�OM��ٹ��(��#���N/ڼ�KV����|�D��䓭�5��
(���	-��zm�
�)������,59pUη��F��� �N�N���}�Q/S�*�0}�)o?$�sX�0-mRם�ޠ�S�;2�^߫�͵pW%��͊8#��0������Mǈ�e�,r���dH�9���u�,�-�y��+bN�8�+Tl5R�C�Q��v8�fP�?{�WSG{���q��#�y$0^�?*�UmΉ�FM�q�?�l��}T ���]��a!��Z@������Cü��<X�������7�^���,�7�`��y�����\N���{z�5��r��i7�Cygō`������/Q�`y���7r/z7��b��q��;n)�d,�1��1����@f���6��$g�.��@�h��0F��`��]D��ʍx�Cae�7���H�O���{������N+��%?5���y*w�l�n�6���-*4�1Ig�w2]��?]?;�3��9�:8�%^.��pxv5��H���
��i�E�;�����X�.��$�>��|x�=\w)��Ap*i7O��≣D��D�jI�/��0%����w_��E�3�
*D��Ms���ˎ�m���2��'�TK�=��]��B��?`�ȗq���	���W�n�|Dk���
��"xG[��"s9  a]nQ�e5���ӳ��Nn��9;����F�+��gΙ� ��ő��cqʁ~��/���ǝ�2��O�b~�$�� ��������V,��Β��V\W�49] ��ZY�M�ͪ�P&�����3���oNʶk�I'y�h3����{���TU�l	^w���X޿�s�.�-��+(P�'a@L�b���1��(Ւ������A����H�O��6�O`	FO\�Ȯ�����>Ҧ���M����q(v�C�?��T���(��E�Y�j)(�j�:�����M��T˴-�t~�g6�JJ��}$�u�X%<�N�j2{�,�~�VgXTn؊����r	�1mR0Un����M'N:k��%P0rM#�B,���3�\e��죒��o���}�����7��*ֽ�W�����^߉�n���z��_�Ͱ��N�Ӓw���D.��J<G�_>>�Z��顾\n��Іr�x �<=��,@NK���M(C�w:]�Y�ϴ��)�"��Fʦ�|`��T��NCTyV��Ğ�?ۜ��#kZ��	`�""�ߞN�ͤ�AފX�),���ù5K�H�VƠ�:��k�Ell/�T�+�-�.d<���ͥ��Cd�7*l�_H��l�ڃDQ�vH�	z�_��� A�Kr���qV�`C�t�'>�m�����j�%�=h�y<���#<J-z�_��g���q�J�٠�<�)<w!�?�Kw+0��1yT:�I�r&��_7L�
H������I��c�ٍ�1��]�����.�Vx|^��RِG0%�R���""�C
�l;�L~�s�����ֈ�k`ra ލ,觝gG�R�8���|��E���̾G:�m����"/�;x���^�#Y������5;c�������|7��Lؐ�.����gk�F�
���g�:��>F^}�gQf�v�]��k��8�/����߂�����Z��.H����Eļ�|D,[��-�|�
S-P��t=�D�/���_.��`���7	Aw�)웨��ʵ�2�ԯL�'�.�X����_;C�=a�z(�P�
3Ƶ����}��Z��!�m&�H�n/R����TA�>�q�\5��z)���n ��F"���>`��{���)������.���&K���3����l*��d��O�p���4��Pߵ��N��f�Ԉ���f��������^�Uة�"��_ІH�T2:���;�7�EEh3b��@������Ġ��7x�~mR������'�ȷ88��AK$�o6�\iM@n�ݓU���ʭ����b��ĩ���`7����b� tJΚ�`�m�|'$��F��5�4�E�,��biw%��k��O��mz,�EN�j��1a�Ƶ�O�_t峃�%Rs�/ˣ�@ѳ14�Q�loh�٘r��Z8��{���-�\\��-#���ԐI���bX�s5؋q�g�e�"܀�~m��T1q���f�y)P����5X�d���I�]��a3�8�c��[��.��T���uS���}X��+��5@�F{.�0dD�.�go� ���%�2�W��^
6m>9X�SR�r*�E� �0������T�QK����]=��ޮ�)����p����Э&�� �����͔�x���yTQ����q�yT�q��vcI�)5�-_���/�h48´��l�C������$AX@[�}Rʐ*`C�π�u9u��[����Σ�H�cw�X@�r�;4ɟ���Eg����-\������!HZ��XCpə�ɚ��E{���ݫ�3�d|�ֽ��~/������X=��7�{�wJ]�gC�Y�ݴ]a����e�4��ފe�7QDn����߫f�w_lK=$+-�.�'�'ؒ�Ks������
ay�L=�1)ٳ�S襪���y�7y������3�"g���V�䆙�P.���YE��8=�\r@2�W�R�?l��N�P[IۑB$h�s���Xi [C�<�ڳ /~�,� �d�"�b�8�2""U���k��'���u�'5�毜�	֑𿅈��o����1���)=�x0�6�b^�{�����,ғJ�n�W�Y�X��>�p�U���|��3{:$bz��{ჴ�x����e�smZ i���t1���4�ʵ�*���i���<���2mI�߿���˿U۩���1m\��;!�.sN������k�g�� @�}�P�������?Y�|�r��u���_�of�&%�F�5|�����l�3D+�o��0���L�ǟY�1MZ8��������(�`}a=s��q��θ�� �>��ģ��bWé�ŉF"�>��|��M���K�җ��92��
f��#Y��Q�?�L�"�6p�D4�8V��y��2�Jn}x��t&�f��7;p�$,I+�x��IK�e,{)�:�z�6\@��OGs��K�2i���}�:M��G�]���u��Nb����;��! ���q� ���u���'���#d��]C���'|���y.dv�Rc03M6<�j����J�'���l�]J�o�a�!g^.я٬��\P�jz���=�Cn�^CԾ����3����O�V$F���&�F��фѴ�(�x'�����H���jHd��k�ҕ}�TO�t�L6�A
F��61S��2{�Ն��R,Wk���DM?%�#�"e
�X\1Y\�Xc��ټ�|���e�m�����}}����H���Z�ӑւ _Ѫb��N���v��C��_����
���S4ݠ��Ft�'��nG�����:e�;]I��K�ce��(e��Q�7������l~���#��ʨ8���>���qS�����G�ab)�1X�^G/&`pJy�9�Nr�zߡ�4 ?Մ^r'�w�L�D0����8U�M��g?u���U�#�c�cJMU����[&�9ON�*+.  .'���!Dĝ��f���&&�K�!��O��F�9HoQ����{^M��������;/%!�)�t���^�������n���DZ@�A��x�������p��=g�ךkνϙW�+w�t�i���گ_�A:�_���ˊ꼿K����3I�W|U�8�x��8}�#��eB46(����
}�k���U
��ţ�5@O�/M̝c@���Q��f�ܐزf�}y���*�.����gy��׿M�h�d�%�-���W⨛2D���P�?�J����v�.G'{ps�w�r�T.�x��,�2%T�w��(�yP̐�U3�c7ޚ�Z0WH<�xA~Ƃ���y� �A�l'D����'�3�dd��?ѼyGM%C{H�1��TN딷�]��2�*f�*8J�5$�fS5e�:��a}g��}���Ҍ*{􆉍��h���wMA����k�WM��~����.	�����uyH�L�0���'���p�~���q�2��%�.�*���GUT�a)	�$�>��#\�j���S1%Z��3q�P@V��DH����~�����|��+xo�����/��H�kY��\�Qugqx8)�^Fg�ٱ��N�%T�6Z<0����!�O�pb ��w�x�*�f�Z�9&��+k�="󓭬�duy�b�7�9�!��Z�* �*F���[|���<ωy����י��{?f��'���o��'w�(t|hJ�{��S��H�܇HW�O�E��:8I�b�@��!��t x�C�%�%��X)�W���*z��U#�|-�sV���h�yo+�'�����?V*���d��������m{5J���GA���r�Fa�{,U�S���6�t)�(�i��&h$���@��!$�i�a���)�샓�I���'U

t�<\e	�m�^�	�}�#m�u|i�ѭa�qM ��虻�q�Vu���a��B~�
{�fш�2�����ԣ{�Z���p5G��n(��/]�#����ۗ�n��I�[�=֣���L�^{���9Pڰg�k�aOHu���
O�E��X�C����U��Z��s�;�9�a�<H)c��mY��3|
e�.�I�`W4�tx�b�F���s�8W=;�c��r���&�^�}x�sa"]�`�aR�{���x��y��_������1�H�Y{]��侓/�����OF~9�i^�^��kLLR�7ɴu�n�?�;�B��T���r�i	�#�G�&�+ :�m)\�2��	H��5��C�TB+r|�|��蕆�(TB��|<���Ս���`���!c �ߛ�V��֬���5/61c�e������N.nPM?��N����X�+�DH�8�	�$�����-���l�}�8Hs�\��f�7}:ǠW�������41~	�"��}}�AB�3��`�X��@�:Ф�m7����,B���HK)ưê���$�Z �"�@x;��jۆ�|C����)B�zKa/���������s>�ڼ��_pS>D��Y��������%cnҾ.˔����!�2��-^�T��G��ї�A�H���n}����V�	��RMp�J��܍�d5�?�������?�����HN�-�[6���R�]wç����#8������]3�d��^?V]��|`QM`��RE)� ����l�[Ѻ��6<��&J�2���P���/Yc���sO�Ψ�P�	LF��I@Rq�\���#���H�0����c��Y[i�e�F����=�8� ����ٸ�m�Q�&�(�.ӈ�],�Z?����r��`�B� �BI+-�ZS{����>v�3���&h\��J��M ��0-ځG���Y7�u�ö:"l#��BTe�0��ոQ��@�?����z~QL	e(��v6t;ƫM��"0����T�Zƨ��5��;���`�kD������v	�;��x$�؋�Q��NeO;�n��QO����1���
o�64� ���!��o���td
�B����,�vn5�ވ';�`�(�D)�h-�+h�l�$]x�$@Z��!I��F�3_�iѾ3 p=�G%꽷� �A7X�k�9\x����=���[D�Fv�����/�c/�D���p�"����lj_�r>�,��]���#���UN�8���:9!��,�~DO�ㄽ���8;����
y}�����T�3�X/�b����[��/��b�]'�^��{�P�I�~����g#����դ�L�[χ ��[���_��b�ݒ�A
�⑭_�O���r聾�����&��fk�K��t\�����+�����6E��P�0�`�b���i�����-,���)���ϔ�o�ߡ�W�f�8
<yu����m��+;.����fO���N����*2D�'`����ޡpVz��Q�Z�U�w���y��mسӖ �5��[��C>�����1�H�۠�/R�A<j@@M�����d�F�C͇��i �Ko�C��䓤�{ߺT�W(>��g�T�,r���?�՘��SoH�imC�`i�
���P��m'��n���򪸸s�Y�MW���!q<�a�w>��m|�t���@kp���/b�d��xYOŇ;��_��$[
{���zcWwÇ ]Q� ���g�\�Ez�ls寵�s ��\v�a{/�Kr�/wL(�r�f4���+=ع���3��O�N2�f�����,��g�A��.b����w/�5�_6pWD{��--�1�em���q?�ւљ:j@� �m����!�8��y:oa��+��|�(�О�C���K�|�ZdS�Q����>dU��ʻ���0��T��L�X�ț����f?yB�-5?E�F�$�nWI �S�6�s�}Z"oH��3ym�hi��=`�v�Hlj9�K�K��1�W��k�y��*D^}%�2�
��� ���O�H�i�������p�=r+G��B�V�a&�HF�����>ȸ��9��){!=*^y����[��
Gt9��|�����n��w�K�9*��;�4Qљ��
 y���&<@f��0Hz�MtF���3��D��p�?�X�Wq��þ�F����g����E�Y2��GҘĆ��嗅3���~$����������ޫ-4nX݈L�P��R��(|%�2�Bs�R8���p��mq�R���7X������B� ���b���7�-�/#"�$��.cW%{��	$��lf�0���y��h��P�|c��C���h��I�{�3�y�vV�~�&��ݻ��CȔ"/�\��� �m�|Bc���$�.��z����?�Fw�
�ۯp�4~:�1�@�c^m��5���(7��2�_G����jH
T˫e��g����?1����{T���/S�B:�8ѻ��W�V����t��Xe��m�����̴��^8���4*4���v�E�[�R6�c����~,�k�Q�ۗl\� ��y��pX��T��]��`���.>Q�H�`�e����6)X�uQ�o��0 �fc�ƭ��J �|��pk^Ϛ�`6?i�i00#S���00��pg�u3�~�~fv�����V�I��b�}4Ѕ�p}+��2�o�d�޸�s������W�q PSc+�#Y�iܻz��w�O�V��d�d"�2�G��L��j)>/��6X��hϝ�(�R{�|�������#%�Of8=c#���}X�ضx�a�<�� �yY{	z����~�k�� ���|�m��[����r��G0eb�ޤ�+���H��Bd3� >��9�X:�L�Ӛ�R��x�Xd�y��c�N�U.%*C$!����?��W�ဎ���$�c7 Z��Uw�Q4��р��q�qo=:Vq(/�,h�9)�X�S>�B��J�[C_��fH�h3+���-h�i��ړ���C��m:��Ō�����M+�6b��49�L3����sF/6I�PǸ�e� �-��G�r���&9��*)�>;��	@���[��򋈮�}�; 5�m9���ä1�&��:��a���V��8�;|U�h���78�ގ�X�B�����=T����p���~W�jߩ�:x�}��������JɃv��%�97�^e���������70ۣ��J���n@���1���qD�&���'�#��r��S����ti�A`�a5@j�%\���*��Z�D�I�7W�(b���$d8�e�L�Aݨ*LK�0^Ln�K�nL��-W�����a"�Đ����/G�ʬ����"εJ��ݳS^� ġ��H�)�(Q�Փള���Ȅ�"�����ٶ��5�B�e�M�3��s��q�7�`਌��e����J�MA*~�B�F���=�f��k�<�ܵ��?��n�gM��_�.e��$)u������NF��.Gt蹰1U��.Ӄ��o.m0
�dt�#	�4I���B@�6]�q��*��+Ԩ�x�&Vf���;�����(c�=����ܦ ]�F�����x�ѴM�0�4�S�>[�U4�[ nm��v�!F��X�3y��-ǔϑu�z�h��J�ϼ�� �)I	%m#C�I~�z�C"�Ҏ�����1_��'��N�T>������4:cI�ڡ�Z�m��Uͥdl��Y��X$O~��^/�-�.����{��Ǡ�n�����{wFL@Z_��c� Qb  [2Wo}�呶���L���W��-�!� �V"�uR�2�����g><��	p�)�*G�'�ad<��o�iK�� �Ľ��K�_{�2eLi�TV��?�y�����$�D�<�.����Vf�����H#�o�9Y���\��L��״�]
Ue�^�":-g����,z�kuq����6|�;N�:3��")�/��C�4�� �Jfڮ�;i�����oy^"���&�y�� �'�Q��+vI#u��_��S��k��ʮ�d?zS7��+
�Yj+ĳ�\�� �`�l���y�2����,� �	���h����vƞrB�0k���������^�
���I� y�C�(����J}ػ�J��8?\ �n÷*S�i�P!�S_��� ��vj�O��q��$i� ��=��JM�z�	�.�H5��>���I���R�U-Wh��[%�AP�Uw]=����"�߉�P����Ͼ��É�}�����w���*<�-pOJm���LW��
��u�v�T!QkE�rLԀ'�����9���ѵ�A�C��0�Cง{����Nn!,�2�c��I�n���R}����Q���\��4����ѧ���m�Ǖ�9�h��z^g��w�=��J�E�;�${)�!�Z�u����4fbB}6g�z�N���g��6��q"�t��@1���biB�a/~vg:�L�Dk�L����r�4	�i9�R�8�5������<�6úC���+���d�C�=Q�9�����s}���}-�Sk��s<j��`��Z��TY$T3s���`�t�+eנ���*�>d*�r
��8���G߄/�Q�up?���ely�ŋŧ��$q�xȀ�8�&��l>sI/��v��|��@��G�m�!D��b��a����a���jJ�N���φ�K췭��|�=�YQ����[䷓/�9uk�Ϟ-�=Cz�����?+�����]�w�XV5��o���r�2���jR�oF,�L�I��X=n����͢���s��`����n2�4�qE�(1xAm�!��2�{N��eoF�	K`�2����pF���ّ��������>�lDH=�f��p+�X��'�W�(F٪G���{L���e\����5�v�P�g��k�:��~[�9y���w�V�����3�����R*�&�br$~���U��x����,���'��떨Ҵ@���DH�h��#~�ye��T��W���^�xeĩ��W'�$䱡R��3H�LY`�hI��}v�"}���5��;N�1ƞ=������d�H�9�R�F]�!��x�5ܯx� ߎ[f� 14��'��'����]��Z��K�%,����$�ڔĮ'�xNmGE{n���:f��Ag')=�L-�U`c �{3�V�;]I�K�ag��>�a6��b:�Cb�x#rC�x�I�hnIV�Ͷ�B¬Ҷ�lz��z��%x
�_&V��!嵎pF�E��5
�$$1]q������!}}��ħ��S�S-��v��j��]ܴ�?^��RǴ�+��5�h��i3H@���	�,~ML���@+���xhRWz��C�)a�f�j�zu>"[Ii��!�6~�}#\!�*�g����p��v����1��6�� hn^{%�S��У��R���
��l��W����"Ǻgy����^�)x����nf���s;ː9Tw�A0������޶��EY&_o�O�PӁeX�loϤ��׾k����*!6Kf�[!�]��fQց<;уdU�fD��E7'7+�����ܤr����ͣ�zCU�))x�fKиue��$�jC�)!$_���ȇ��%�S�%t�}�#:u4v�M�d)���>&
�ތ%ݩ��[r5����Aژ��;�(!� V5|.��$(�������h ���_�s�ǈ|Φ	e4�����?�Ed_�6֐|�j����Z���c�ZV�����ot=��q�ב��P/�DO&ח��UBa���镐�Ѡ;��:a!˭�:�6+䥏���Џ�ļg�h�A�>������.*�6n.F}sb�}�E���L0s]OU+3+}H�2n?��;�Z�M~���4� ����,�}%ߙ�������5�Y�ѐ�B�c=R����<R��;k�lف���!��#�#�Z�~�C:���ӂ�܊R<D���YqBn#���o0b-]���'g�ӡDF�ML,/}�f�w(�}�h�fg�Z�����<���T�{���6����M�� ��U8�|ȷZ��È��9͓~�֭��i{*���HiɑT:��6��k�[�������X��<��b_�u�:Zυ��v��:��(�&�Q�$V>���Zf�gav̟kk�f�!?\U��E�)�\�)<C��2���U^X*g�X�͋���Z�5Ri�x��\RR�?
zs�s͆d^տ=��q��w:��E�S����A|r�YJ�xU���,�SJ<���ղDe��t������*�$D�i ���:2F�E�L����IX@�Cu`Q.{��
yѷ�ݓ�}�;��%ܡPhn��^����Bfs��>ȳ�r	B���4	̴'j:h����XSq��������Bf�Ӵ��5��������Ġ��sTD�[��O�o�z�OJb�;��e&*�Ӛi5���L��ב�z)�n�,F�):Ac����8_�i��������v�/��1�jD��k�W����P%!�$�ҋ�]j���M��]��Q��7�:KI��o��T����A�o�kl��3|%��Ǜ��K���,(�n���NGvub6d]ʭ���&ҽ'.�]N��� �ly�X鵮K��v㊰�.^�b}!Ǎ�L���=]�0��ZA����ʶ�fC[�E�m�}���-߿�����l��T�ӛXî$o�/��sm�pc�TyJ��(pR�D��H�,�F�r��������(�Qb�s3�XÈ�����J7��X��$�-%FQq4o/�~8+P����R<�\%����p4�N��`�b�T2�TR�.2{��tFodh�..�c�Q�?��<�NX;z�9��B�YV�JN��$��c��c �u�7h�xQ]^\<��¨8�T�����Hu��DG�o�nDT|��nYߨ�#�k#"r�8�XΗ�b�	A���ڂG��W���TtL��jǪk������e)2l�d�͢���VH�����[�c�\�99�dв�z��62A3�E�
Z�^��ă�5��I��I	��D�J���O�����V�j�s��J�NnudT�PS��8��aE��̜2h�3B�m��n���i��TK��ᦑ2�E���e�H\��CУz��Iu�~}ʺ�^��O�Y��{'��a�L<�<�%ͷ�������gM�U g=vi�d�'��7&�֋�Ȧ�|,�4��O�3=�el�M+ʼWZE"��]u,���t��o�%�׽:�,y�(�v9 �qHēN�P��(�eŽ��Y�a�.�Rr7��'�v�uZ_q}�����ઔh2�<E����׏���i������@�Ġ����!n��1j͐�q��B�J���O����5�w�z�ؗu��4/��"����߲�	�$�fױo�xg5�-��2��6���<����F��1=�6c-9��Ϟy�G��U���Jd&Y5d��	FBXa+:�S~o��q �yT�Ή벎B���x~V|`�V!����}��wh��������E2�Oe�؀���������)*"l��n�:�_D$N��ԭ\��5�(���+���$Dt�q��F�.i�T�H�����C�h�5���eF������!/Ny�f?�O���Z�d-v�D�|R�-�ui����$X��?��9��6�£o��q�f��k�����s��_�������Q��~y�rƦ���_ekn�S(�};��� �K�SJd��m�6qp�X���DC�2����Ȟ޾�B�)� �}�S����<���n��:D��@A��#��uz�N�{3��Y�"zx{~�b x� o5���a͐Ђ��6�+��5�b=|���r��0r)�h!�B;���lC�r�7���\�d�a�4.���t��t�3?r�7�g��P��I���עaʶQ�앖��(Y���qx
!�����
���� D��0�°اYZ��1�`=���4!�c�H�Ur�V��n�tu`�g��'��|�uQ�|��%������l��Iu���kn���1��~��L|k�� HK�Fv�ԗ_N-��GYR�J�_TN�Y3`AU[=�-�@��ٻ�?�P�B`*�������!�!�C#ا,��=G.�*+�5$c�^����
�T5a�~�I�����(�����8�Q#��#�Pqwǧ)Z����o���M��{����aư��Wy�s助��tQb>[���1�a1袓��0�᎒��q˛@^�~�1{�2���a��8���n�R�K�	�n� �?�D	d`�����������p�Y�g W��
p�u�nm^&�{�� ��|#��@�T��!W�=[��Yxۼo�E�6J�i��j��oy��a�֡��`T�-襝�G{���H	�9���%D\�g-)�H�����D5`�+���m#ݯ¨�����
�?�����Ũ5Vf��2��[��R>�`bu�S(��g_��O-��~�nz������~E�I����̇�o)_襱�9��~Tvz��zx:�y<�]�����=��t���Ӧ���H~���r(�P1q����ױh3-����?&�/Ɋ�H��s���,���Eb ����OCP�f��p��m2r��#De�̰��&M��2za�	���W�����U�۝Z�8U���Y`����YKn�C�g5E4�_5�8�$��"' ]؎��F�:"�+�N�EE�Q�~m���.;�N�`�`���\����Qx�*6 �|T��=��m�'}?#����X�>I�Xj��,��z�~ha�Sx?XEO��3�����1����
e�``-Dx��U6����	���1b�l�p�q�)2A�&]�F�ڂ̖��Z���8(�;nc��)��d���sd��}�׽j̶����`�p���-Km�Gǟ��%��@]��X��E����5���&

�櫛�l�Xi���������P������"�b��@���N���kG`P/w+4�f��eJ1�K���� M��@���(�2B��Ys-�3L������������ �ٹ⇵{���l�l����:��r�J�� �%9������TCL��0�a�-@%�z�Tn �B	�3��ى����_�=�)�����g?t�K��x�m��.m�V	qc~��X5]����\=A��������ݕW¸���f^����W���]g��@�����{':�<���	ߪׁ��� Ă�h�, ����إ_�e�}܌����U;��U�"��]*���D�NJ�m���Z�'(��ڝ����"X0VM1�b�B�a)�㹄���"�)����6J4��XS��vdt�(W �UH>�5�0S��
��Bhl�Tv���@^��8�vנV�9����������k�	�n���}���J#��E��6�&JX("��Ur3)f��"�d�X������q0�PXXq.eI���٭��EK�iT�h�Rz�a��zB؈�q�������C�;_��O��τR���+��6��]��2�gvA�,�q��AN
??�� �
�L�߈�����}��>�������9��dd��d4	�噱�Fl�w$ˀ�߲iT�)�7Z�hr`�^	����oDG~R�Kv�%C�@D������D�ų���D����t��h����%J�a^x��ZwȮ��?�>�̒���sf��\�#����L�D9��_�����B�p>3ƓVc'�!�Oh̨����gH������E�f�C���G`n��F�6��o\}�$�c\-��5�n(��e.������cvuB;] ����Deq�m\�����o�rɱ<x$���@v��=r�\�����>bPb"s~���5�F��Ƃ��?-j�"�	-�"?��ڇ^������f�_1f7��t�t�����`sl���0;���5�ĳӷZ��}�RT���g��I�E����aJ���1�7!,������vQ�⧘726��
�Ϭй��BԿš���z��Ź����&�­#�\��tK^��?���z���t�N�b�+.��I�h_��o���0��N��"4+Z�3�Tz���G/��@�"�lJ�(Q)��'>���3� ���i��7����7�ˡ�$Y�g����^>3<c��w�y�p|�bj�M |��TKO�Z�w>m@�z��k�8��J��Ba���|���V3��X����$c��lǜ#�#�5�z���I)���v<��?�`�q�����@�7 M�2�S��Zz���T^I;���9 -U̡N��y@���V�#���}�R}50��3� :�D^	���B5�j6.L�T�<��,f�� 9�7�0�U�&��!E�
2�V)~�VpFN.'Z^x��"_��\�g�3
��=���­�{����7l�|<u����x�/�ʌ`G ZI��X�_�<�c��Ѓ�EiN��Y����<p���+#u�9�V�0� |V.�5s�ę�L�w���RΑ���e��r	U��CU��I*���^A܁��F)��1�G�ُc&8}tԟc��$� �� ��1b��Y^����w�@��ƺ���e�� �h�S^� t�Vd��&[����le�(R�H�I?#=υl<Y��
��w�:�D����^nT�n#"���:��:�i~�Ȫ�Ppq4E>��ˣTz�:WF;�l���.�ڻ�H	=�0�ޟ c�-��m���9���"�FeV�y������1����_�VtG��̣����M>K�J�[����= ^��~��k	���(&�"��N���6*q��������JF9���W�uA就��g�L����Z��[�f>�����X�Q��Id��<�&�]�Uz��2�h�=�� ���3d�dTܤ���j�"Z�ͬȜ<
5��tb�0rT(Ɛ\	����FY�lm��x5K^u�� /Qܪ��F�|]�I	'��յ�RC�F��wv��*K�6B�1f(~;ι��E4���	�j'v�M �8)��w��|/`�K�%�L�a��QHS8o�͘j�%��y��y��̂�~ �I2rŨ�K�\�0���7�b�&��Ǉ=��N5q�-k_@y��aH�_��8>C�C�7L�"� ��%ڀ;|J��(�F�W<��P�8���g����CC���4�rؓe�c[<q8��8z�]� l�=�������D����YX�t�8��=M��N���6k�\׈$�.�α\�o�%0aN�ߐ���-^��p������/���5 ����\�~�J%#��E!��5��%L;����
����-,���  К��y��Z����Q:���ʸ+��Ȁ0�3mH��EP�&Q=�p
���dB�pX����,�s���\
�ycN�8YՄ��[��Z�z��䃾y(/�L2�}�O����J�P�d̃�C�ja��GW�|��FD�ն���ɐ��h��Ƃ�	�Ȣ�e�� ��D�������,�H����a���~��z��V��}������z)�=~��Nj����Y:���x.��m�q�|�O��؍?���Ђ*��[�<����!mP������w��v�A�x7V�����$����Z�exm['��Y�A��n���1�Z�D�._Z�tJ|�1�K\���_�}\�a]Y�0��.k:���(��L��GcEN�J�(ϾYยKE�!m�����V<��ׂ>OQ�Si���������&;	�oJ�����J����n��	'g�Er��+z�G}�;�(�W$xx�is7_��8���CJQ[R�'��O��K~-!a}{��L�a�%�͜b��G�	B�a���h����;�\?ˍ�Q/��xc��`I������V���@�nwb��vtU$����DGBm��/U�����M5ղ�o������%h�~��ͩU ��w7��O?��g	y��
b��ʋ� �� ��v�K����E<�̦�Bm��A��9�B-@+vJ�"�Íp9�N�Yn�u��;�x|!������P;NxW�w5'F�3�����7z?�N�F�̐o+�-#F�6L��CuC%龕U�+�)A��{��e�w1)�Ps�j��U�-vSB���Z�w��s��@afk`}F�i�+�i��!ˏg����M$S��RYM �5-m���:oֶ����W�������3���e-2cdԣ��Ϋ�tβ/Y�-�s�ǿ�s���QN�Ħ�=Sr���H}@���}_s���
b,���a%;~��:�Z��c	�|��j�m��PT�؈��'�5�x�, ��UUҢ���!>�f������[ �Pw n�J���է��\-,k�F�����8�[�A����<���v!�oaPuMCR�]��~ɎR����7��!|�拱T9չ���/�e��[9��J���U��.wm�֢�bj<��^p?��X1\Hy0w�"�sv�x��
�	�{�/_-���E�����=���s����������0�9���t���D����˵<��XA�&*%U�G1\2����1~��.���K�B��d���!]� =C�t���%O��y��V����*�q�S �6�h"�)��_����ld؀9t�*B�I�ه|�?I�w+���*�^1]�!�ͬ��N�.g4ׅ�i��\���3����d��J�D�5�7zP�Z�+d�%���+��i0�}�V��7�oz����P�(�dLG(x�l%$V���k��]��k�t�#!�� 7�y@?P��#	v��7\� �� �
���N7b�C[m��ڧ;�+�,�;�}���j�m����\��lϸ��{O����Q�@��g�'Ip:߄O��k�}� <�Uf@i	v�l/��t&Yˈ��B�]��n��b`�X$m�a��o*�-� �k�z�U�Pۙ�P��믻��s`M㑮۲/�q���д<�8���U�¢x��6����{�P���'�kc7�Q�տ�( ��_%���N��;��r����T%�X]y�و8�=P�rD��������� U9��Eba�&َ {�2��E��<A{�����p��'o�Mj��^5��L�B,�����ﲆ���WP8��D+鏮.���=�t��v��O1��>�z�Μ�|����+�~���B���*�"�=x�wΉb��%**�Vq]60PP/�F�(U(��I������Q��0���0G����^�9�7�'��G�k��Uyx:ldA��~P�Zw�
b���.���릥����Sǟ��UG�ZC�!�[S���h6"��������1�n:�����ߙ<��8j�u�s�`�������g��N�+A�0r�ru��ԙP���5毱��	���*��}b�XB������r����⵫���,��Yx��`6�`S�]�6�~[��E;��=Tr��!�v���-���Q��U1`p�@�o���CL�h��3<0��V '���<�,�Yn�U��ڲp&D�h�!�	t� L)��s���D����O�y%��H4`Qii�f���]͒� qc��y��{ԍg	 ׵�}� ����~��Zz�}e_�{D܅7A\��G'.��|��S� y�O��fc�O�窣���
�����*uXU��12���JU��<��'�{*�=�9�\/�I��+���F/�B`��'�r��(<e�Jc���.N&�w���P6���S����ʀgA�$�����O�����Qǃ���� �rV��@c�Pum��@0ё.��5�P����XOƒ�9����¶\�y���JL��6?�6Y�2��xU����q@U�
�<G��e����}��!�3�xܐ���.�^�Dgg[I(����"���tj5�s�QY�y�����NXx��!�:�g,���%˽�5%�!���->�s��D�U���x�Y 'l��o=+U����n���<�}�i���v��4�ߜ���U �����X���U4�n���F��7ћ`E��x�$�?>����D�_/r��1{�B͍��%���X
Y���Ŀ�H���-�"،�N�ɿY`����i=8>��{��%��&9nod6�g	���(�%y�?���߾�G��ױ�1�8K�'F��q����";ӺYA��􀵠�T���f��Ә�a���X��T�e��
����Г`�ֱ�qf�P���^�����KЩ+^����7���h�m�䂵�(Z��"�}bP�w��!��x����ςP���i��W��	�����#�;&b���cj0��q��nX\Y_#��%N�2���EY���$n"�6qF�1���=�4���u��$QTf�(�_( O�8�KGj�+!�OQ=�/(�x�9d� ��q�k1�e�����e��PĽ�YyI�+w@N��8A�:�:F6{sl��!��aZ�g��[�5^t��|���DU�AV�@o��cJd\�}�Ϥ�� +%"}�#q�7�un�, CD �d���d���@O���(+��$g�0#��J\�ղ�]5'�S�c���\G[.��f��dD<��1v�ߐ�m%`П�W����؁�����߂�������M/�A("����V�)�)@r�k��&�C|���bCa;^�X��NF��<��1��/0�y�Zs���C��7����2����}���or)82��~����p�n��$�����)8c_2겦��+�����Qks��r�
�e�bz�h$��������#�6�6�k�X9m�3���m^�_���}�{�	^,?_��"󡒴�&�������3��vv��N"#��D��=eƍK�8��y�c�-���
I ;���z�O��}�~�87z
_� )̏��D+:�D�5\C0�\���~:jc��t����,jR��[�����g������o���P�p.`��A�`[Q����L�];�F��N�kITA�ʌ`�����,��wEt���F�r���AO-���úݰ*/��l�޸�t�"̐J�F���>G���gY9�J��6:\?�"7�־9����#�	�/���Q�]�xn�g���>��oY���ԯ�~��E��U���_;렱�|?4^�";c�8�+�*������}�7RYnh����X��IK�A�S�Zx�ߦ{�of�1Iz�q/?�������|��� ^q]�N5�� T�i���G��Z��a���&*_�v���%vkg�I�e�`�2#*uē̺s?�k�lқ���^�
���'c͹!	��6�Uj�����C���V�4��aF�9[�[c�d}P$��؝��f�r�2��D5�Y��� ��=�(�E���[�=ڗI��B��4������o��T�J�bKX4���(2�/W�D��g�1�!�K�|v�19U'���0gx.葳Ύ���Y�M0�^�Q���9�/���)�,yhC���Q�b`nN@��z	�L`����cJZ���ҝtᢤ�}l�S'pkBH�˭"h��ԿX��hط�X�c��j=���iٻf��9��4����H,�"�<u��/�^v$/L9#UN�(��Әn�=����(S���u�:��5[�[����ED,���u�(Z���=�w�?�u��o�QG�.����� ښOq�r��=?�\���oE�����6��\.|㬗оoiJ��qtKJ���n�����>��v-ը�7�ʭ��& 8"q�.�Yv;��޷�'�cv4.�R��F�|�$��=���c�k�tb�l;K�v�cWP�f��m�����<�q"�1ӳR�N�dh	�^��l+��"4Iu$���HJN��{�������9�������`b��kW��<c�����[D����O�D��x�qb�����~��/(��p\�"KF��
�#���0X^�y�h6�Dm��u��&�:��D)OF
�7�<>�W ǌT�%��b�c��Ѧ�Y�7q�r�y�MzG
����g�mS�	��[W�ɏ�6㡘k���h5mN��jᓘ����I�\̗���w�9��f�
kf�����,�)�XV���h.یm�c5��(cnb��J�����Ig����g5.�rdX#���ǔ��"�\�1^gC��ȠeZ�>�aSz���v�	W�v+)��d�=W�}{Hz�Ӎ���c�7�[�p������IC��.	��+�J��$��L�(���.�ܔ/�xF�ف5ԫ��@���vP9��O���&ECJ@-���Dhr�Rp1�ɵc�x�#axjv�1�U1Ty��H��3'��a�+ت��vi��n������[���i��K�[�)��ֻ6�������nu����c�5au��D�񨂘�i�r���h�ދ��a6��ž�[~؎=f%��R$���Y���ߠ�d�$��Z��/�ԆQ('	&�x�g9����H�N�t�w��-8���;i:LNFE�(��Q"���n<8�s7��=H���CMU�a�G�C�g��f��c��?j9\�ܦ[O��áɭ숢��b��}�y�Ѓ#�Yb��0v�M�?Y��<bAC��Äe��Xo�ߎ3�5�W�a�@�=,�����@ÍE-6��˨�����1�x�|@9V�-�R�������cK/�?m����P���������͎ ϊ��/[����Q���Ic�˾�@j�w]#�1�T�	�6"/�
���Lc��l֨��t�m�sTN!�,�T�B� ���Mb|w��'�߀+����4���ۿ�<||�~�`��^Q�$��eH����q"��W�OH�{lԐk�ڊs�'�Z��e���e]�u�1[Z3�����@���M����5ሽ��B����#��[A�ٻ�*�0����e����Ъ.-K8�_>�JK�y=��R����x�5!C+���Ҩ%�`��%ߛ��	�]�H�c�j��M�).�eD�TM�M�~�M��R��i6|�^���hͱ�Y�?���<V�,�)8̐<̛��'�u�~��7@��?��]��o֝b���g�J�^7�������rEy�y`	���E){�Q-��WM}e�w��/a�"XG=�c2@p �e�\p�I�K=�ot@�M��R����щ	����<A�dba�m5"ͪ��Ă��[l6!��gz������E�Jd�PŤ\�/�BO��l��!s��E�� ��X筀�-�K�Tk2K�'d�J�#k&���DdT)����#i|��U��<'M�-�Dm �pb�7��uBD��uӥ�����N�A
�f�|��1&C�B�@� )�g��m�@mQ�S<�'휭��pSH�(�'h{s>��w�uB��Aq�-�fX��L�Z����Ev��8;����1���ڷ����_ ���//��kq�"�����uf3Xj�k���n�վ7mv墳OZ����BtՐ��3P�C�r�p;:Q��9���N=� �G��ƪ�؂\�G$M����1�1[�[I��,��q�Ch���b�7K��/�Pr���=��u��3_�W��Mke�_xVpc(5J��T�����Hro<8�Gt�&Z\��a�Z��~��1��g�ϽH"=s���u��<�%�A_�xG>M��P�M���*"!�'�uL߈�	ջnL(p ���������E���:M�ɲëI1N%��� �� �����-sn��m���:�mCQgM�9����i���w�S'M�ۇtv��)kr�"iئ��A�_QW�����kB~�x�o�5�	��fs2WcS����3w��)&��1�Yc ֥�P~�MiRC�m��$�^��h�_8�f_��7=���S6f*/�M-�/�� g"ף��!���Go�G'*8�C��+�/�	��Y��{V\��|�� sXOB��W����R�g�=��Ы�8sV��������c4�����u�Rz|\�6۽1�K2:n�R�3@��5��J&m��d�{.�tc���aI�V��8��2Է���g����
���U�^��`=u��Q�#�(1�G�1w��xS�5��ڪu���x��@��\�(>8�I81�t�mm;������ւ�ߣWK1.���um�[��9��һ���LD.�j�b����C�"�{"���a�cJ�7�8�د�����a}�#�y�y��j���F��Tؗ���Vw���Ob���k�?�?�l�̵��-l�ya�h��q�$���ob�����zg�1X��K
�4�9������ï�͞.��|�O;(09K���5L]N/���E���R=�i�=����b�Dk�w�]���&ϙ���ޓܛ.ƺ;��6ke����)�M� �m#/ZZN�W�pc_��S`�'���C�<�"�q����6�N-%Ȱ���N�K(߇��Tt4���9ׅ#]"&�/�n����گr�)�me�aR�=��.4���>,|i$P<&��)�����T�py��[���o8�!ܾ��?����ݽ3J��B��}�G�!~Kk��M� kN*���y(؎b<�����8!a���'�>9��]
��k����s~���w�!.������t�������Tc~[F�j����L4�˾��� d�����	�m� v��z�Y�\�vb�<a��,�ka�o�m&+3�c'�G"��b�1��^�f'�����8�$�������DډO�Æ?3�������ٗ네bE��y��_P���<��(<��t������v���6�೨fШi�{��ӌ�8�	�,�����Z}<O�ko��r��4�w�+�L:vE�W�kmT��������v�ߐ�Y��3���>�xS5��]R]t ƺ�E�@�ߦ��ҭz��$	'8ѻ��?<�N=�^P%zG��L>���D��k���&!��sU9P���B���* ��IT��ي��$�F�+\�F�S�"YLaV�aR�MK��۶�k�!H�[R|��&
�ƶ�g
��CI-Hx,&��FM
ǂW^^���u+�ݾ_s�V[e��kbf
⁒��Q�ݳ���Q޻D�Ql]��x����k�I��$� �R��Ɉ��aj�?�ef(������>����j}IX�0�U{�^���[���wWy�������m�z���F/�_s#zh%喪|�i��<s�#zGd�P^����	!8�ι���n�q[Ά��Xe[;0����m�3�� ;Sm�j�N������y���iEQ���~?��U^�� �M�;�����f]й�l�鿾ȹ�2�
�9�h[�C��qQ̇(1EE��J4��}�����~A��f#�O2ң�L�Jz7q�P�i�ݪg���?�\ʮkt���7��1��,�m�أ�j_�>�F$o%�B��p-#�6+b0@��dTo�Gi�ܾ�Ʈ*5�X�I��z��=<ᕘ�Y�Rg��M��Ѭ���Z|��4�p�����9�L/�p�(	�����rit:�N�j���$c�-�ݱ�A���NLs.E�L#>z2���@�jHf��q�*\���52��p�\��e��N_G�X�s��O��N;lo����T�X�m'�/�{�EZ�&���"P��&�F���X|�8�z�U�K~a4j�C�o&ܗH`��6�W��KG�O�������H�B}�Ex|د ,�0h��g<�Yi1�lV�h��"P��&f��I��V4>/�J��x��E�d��ܘ?�ru28_>���+38�jw��Y9<\�cǌ�sab�eLL�ť���PH�9f�ڊv2e��v�ya�ʬ^Iy6���JC�e�1:t�7� m�`�����L^�8|*k8C��C~��_0��b���e�{%��	RQ��6���)"�3u��	���0�!XF�*�U��~�ޮ�~�G�H�j�%"8�k��ۨ��Y{���þ�h�cƍ�� ��\V���7���Y;���o��UUu�e���s�\W��m>;@��>�[��iO�q)��SG��gO>Iw.���YYqU"?v^�aXF�v,�I���ކ����N@�?m4��%ſGj���/n�M?��4l5p�͊�����o��-���EA�xw}�Z~n��e��7��'��5NSJV�ų���0��q��B��x`˭"��3����	�6���6S��LS�7�?�S�Ҽ+�.�9���OP�3z�e��u���</�����ϷTh�mɕc��I��QY��Ȼ�Oa�ޚ�;f�� �-<W��ˉ������#9���c��5��sST $�,�ѱ�S���e��'ZB�q�Ng��@��aZ^X��p����U#��_�2�Jc�Y��Ӣ�bM�t{��	}H"V��@�{4z!�(5���.�VDa��	�@@%2��|63��y�LE<\�ݣ�Z�Ce�۱*v�P�W4��V�jpSs�7_�u��[��p_J.�Z�3Q�q:�At�[��Th�c�pRL?��Y]��:I ǦDr=7֌�#g�ܰ�9B\���}`���Q�> ]�������fmZ�p��a`ptӤyڥF��4Ϥ�H%����5&V�?�<x�h�r��K55��1&�t�T<��\��SNC�� ��W�`~�e^7����7a�����R����fjI|�|@r����׎�h���4��k����1���-��a������N�_����"E��ێ��;g\�V7N���ﹻ(*1��,�V���)�а���ᔕ��E�@��O&I/�&,�o�d^�Ӟ�ܖǬ\hu �ǳ[�`Ù�l6) d �:��o� �z��c\�?<x$*s�[�T�Bg.|MԸ��������E Y)��(�b ��!2�>��`��q�gn��G�HA��K����eg߈%,N{�Ǿ���mNR��O��&�%�ts� ܧ�Ж� �&�����2H��>'ƙ�<�H���D�q�sF�9�9(p2�s�M>��Sm}���!�
�!��a��~LҰ��>i7%���v��ră`8����q��f6W��u�x���p���*aj?�˧�.�G	�գ���m�yTI�k�&R��\\��6��2��������Z���I���k5�ZΙ�`���cA�@J^素����P�q��H��Ѵ"��b5����#J�K#��-)�����Ug��r���̀�
x��*�gSw���쁘>�1=:c��;�bX(�>�1�=n�Q�ُ�!�\���p�j����*>����}��m��)�f����5b@[�B�U��o�~�Y�NA����ȌdMd����̓_�V�� ������ �w��Y%��$B��m���`�٪���Tio��Cژ,�u������:���]�וg驥��������^[�nm�G�'5<�H��N�G~�>�_3H^=�Q�v3_6rn^�WץI����� e_����yf���_.�G�`$\b�v0��l��$sn�`\�_5199A�}���i^p4$��B��bM� [*�K���C��ь?a��^�0	m	��V����ur}����zd�Fs<;W�����>��=k����k@�ɔ�U�.�$����>Ņ��N���ٮ�ߗ��`�6�
jo�/r�a�15���1� � >�S[.�'-��x����[��3sM&,<�����'�*�UcU�xP���nH.`�c�}t�V=�o���i��?t}���d���.e#�$a�-6٠�"��G�2�M�]V
�_<�����{؀��Nm*�{��3%3�)`^�p>������/]6
�ed���1�ɧ���a|�
?��(�՛���L�	�'�O���j�6�ǎ�LQ,���Ǣ����6���gReU܇�=}���ѧ^?N���}�����rx�\0sy+���Nm�n���2&Yt��f��[ݩ���47��ş��"lzߟܪ�4��0��[�_>��mj�lOƗ�ь�O���� �e0$F���kR�7����I���t�C���b��趶���A�(f�����Ľ��
qؓ��ŋ�@����ۆHB��s�Gv$h.���MR��5�%Q��`te�LzdrT�Ć']��sT�(U��%%�i.���i�.�G&
���� i��7�n�����`�����6hT�K�պ��r���V��:]�7��4�LY�֡�w���e3�Z��E�w������`�5�_���Z������7��9>��k6< �=k:ֻ�c7ޮ�4ݔ4�ZNTZzJzy���{Z���2v�T*��I�*�*����s����:
+o�s�xp�,�O��cR$¼��E�<R�������3_ -+�ov�(�6��zC��J�v߇~�y�����5�6��PC���p���D?ԡA{E۠��i(�=�_�܉�-�0�|����ߪ��mj��7}`��)��D�����m�����(\tM;�Ƕ�sn+�F��� ��G0��os������?D^�jWa�Giݴ߶������>̤Ӱ��ȣ"*^uE�]z����c�p>�a��prab��3{����'^A,�k����,�詰*!y���;�Ϋ恺Κ^<B}b'�|6��U򘂌��,�y��8 D�F�$H���e�,����ĆP�e]g9O侎����ǰ���lv�	T�b�'P��+b�EP�"���-^���7ƓY��U�.{4���}�g�:�b[�ϞE*���h�͡�ڞ[ߙ��M��_�w�[�/��_���V�ݵ�`�`:�c���{�D�h�at?��ӈ��Zq�ƕ<���Ǐ[_=��#um,6E?x��#�]��6���&����b>M��A'�v��G��c9p� u�Z�Wn�30g$|�{g���������]��=~�D� ��K_��aN A��X�d��L^67���tc�8\vbuv��:ocedpRO#p��FF��خc8� "�c���1�<�m�T�-h�'8�׵�gE����6����C)�5/�SKu�9�&�F�Xӯ�\�ׁ�$��k�1��w1R#0R;.P.'_�=��\�&>&E�ȑ|5b���M[u<�;��h��(�[ˈ�ܑY,&`�ڵb��?�w��Z��a�7Q�-��d������P.*����&hf�8��y�z��E�Crn��#͖%���U;"8+���c9q�w����F��s�͜�]8{X�>t)D��,�A�
�¡��0��j��/��ĔnM��u�@>��X ���fЀ�E������|�d]M[�&s�T/�]'�4���GE8���ϱ�,޵�q�)wϞ�(��^gɪ�<vm3�Cܿ��~B�����P1P '�/��Ջ\�@^�B�k�3�Wq+�^0fx�)��]¼s��\���	SH����u��^(���[�*��a�[���*�ǩϑ�G~�޶C��s�b�S6f�H�������},��:�=�Q$����~9~��q��q��q/�d�R0���;̭�gdU�R�Պq�`�zb�Q[��#!s�=�dގ+p��x�R6���ʺ�Q�}�}iK'tf$����ú�2n%���vB���:Ci���������9��]�_�6��<��g�1��x�k�fk��NEQ6���;�EJC���v���b���1�*��ϓs�D�c����ٳ��r#�9�yӖ����CQ�sؓ�� Z��n9�o�*̠��������t��]<.so�GF:��L{ �=\._U9�]���g���Ha����z�&#X�b��մ�뮨��6��q��H�M���냠2&Ɲ7��<�$�,1���
��o�py5���4˖��#��BP��-t`3��fȂ��˯�4���c�L>P�p������$�@��,�soQ�9�^��iJ�������@@\�a13���ˁ�b4����MY�V(KI�1��P᠊��lq�UD�]������1.�"6I/?R��?�W���$<]��s�1�����m}h��|�~�G�[/���oP� wv|������|�Ì~�r��Q2�a[�'�����%JUO��i��ۼ�4;��}�a�LJ��ʯ́��~Lh���-'�������漑�b�-[݉�j.Ū��]c��'�����G� y=}\�|�fύRk&�`����2�^�u�o�yt�����:P�
��\�����b�ԁ�Tr?�(G%d����2���L�ؾȠ}K�j��^K�IHdi�q:t@�����6�-̒=Ѳ9i}�f�b��rif�;T��j;���ϾoӴ�(�|�0R���VO��,����'N�G���ݜ������`y�_j�vԇ�������EͰ��Z�F���e�UgA��)�p1��H�n���˟)K\k$�N .u'����4p�`ˡzE��T>.��W)�ypa�O���y��^�KQ��\��8��P�-+�y��
I{�fN%�[6q��-��_���|��ޞ�2	?�1Y��BW��@�Xu`�Z�Q��$A��E�n���Y���/5c����gxt�ީ��G}�_��R�-/������<�V��r'5 "�ԛ�z��S7a3>�&��A���'�����F�W�;z�>M��pd9�{��f��1���Y���0-]'$@|��
I:�vv
NX9���E�P�*�Y���7 ��YH�\��"M-����p^��;4���3c#�Vb�� )U��JP.�z�@�Hɯ<氆�ڼ}��Wd���]�X�m�f��t�h,[Ns���/����"� �~�4&�畄-KE[b�c,<�� p{�p�f�sh����'t叄G�a��eN~@m��@�zb�ٝ����c��[��i9���7r���p�'<$ �� b��FЯ��"lh���Å<��w.r�������:[�Fst�N��F���4��<�⦝�|�[�܂y�qu�g^?�&��7ol�{^����R�.���{N�i�?gYi��@�+j=wp,u�l�Ќ)�5I�RGo�5,�->5����?(
0���t��|]"Jt��Ǥ��4r40���a�F}�9>p4�W�#B=C beJ��n�>��B(�
�'LSwI֞��9�"�
�w_����oji���>I?�*Y<���J���(�0r�F���ƞN;([6�B3/�" \�V5��� �bY+Y֏�]�6o��T�ދP%]
�2�@���:��9J�!�|�y��d/�������Ŷ��P���űm���g<_|�>�w#��;	�&��_�4�����5^VFy����xa�tE��1������9��Z�j��&��V�/-h�URV�m8�����������/�c|�2�V�~�����˪E�J-ak��H�A�遜8+e49P�5m����A�����kW9�a��w�*;T����H�zl�q�)�O!ٞ�!�|��<>�d�?.�M
��X3g��/��;����!]'����<{�÷hK>�0|�0^Y�-S�Ȯ_���Z��<E\��=)'�x��i����=!5ytI n�D��N�\���ޱ�K�'p���}�E�uߛ?hB�r�d�<�������;�ȇ��)Û�Z��?�|Fvt�Sj����UEģh�`O^Z���^o�"FV���np���qh�a,�5_���?� �.:^�u�ҧ�	��xʘ�"r���Fn[&k:�W��Jc�*�w����r����{�[�ˋ�������P'�6�tA�5�Q�����*��ȑ�n�ןe�o�w��/g�����o��âQ��u$���[��������r�; j�������W��m'g�p���$\��nx�qQ�����N���p�G�25)�sT(ܬ��1���>�Y#�HM�,E�IM;p�铿!B�������ʁ�� ��
3���!c�¡y�v �"��B�2!Wx�ZcP>�B�x6j=��
����C��o.?�����-Ǟpݜ�����`����5�FD�xeW�g@���:[�f�~Y*�}�/��<�9�9�D�IQ�]�V�������A��� z�z��B���"e�����|�^�G*�����J��B�;��e}�z�=t;ٝ�Ȩ����s��t�,qQ=�_Ǽ9��Y�)��v//Α�D5��Q��Q7މ7<�`����D�T�:h�R��oy(M��d�p
7�b�vC��W���ڋ�Y�f%�"d��3����?��~�M��H*��0��I����
��M��RA�f��������^��ۤv�;v8X�oA�����!Sw��Y�n�^��se}�~������2BwAtݺyO��+$D��aً�E3�w��l'\:ڹ�|��U4-���'VM�v��i����:�Dx���o�Χ���4ӷ�"��Bk�*}O�a��;hPR
���<�f���>��m5�[OV|�՚��}Ri���q��ї&�A�Q�y�o�Mܑ���4Y��!De�Jӿ%�4^����9Li)���(���P����6�l��T7J�T����Zl�+p�=�|IΆF� 2
D��,�Y�� ��)��d��_������m�g��q�uX�[
�f ���6�{�s���ش�8 �☉0��ާ���.�E��� 0�2��ZW�)�+�2�}�ˤD&�Թ�J:�5lP�����������o3<⍤i��u��򙪋� n��nN��&	D	�]�_�\�� ���2p�O=�����c*�t\���ZֿC���\
;�� ��6C_�x�X��h�XxV.���|�q9V�7!�(�.&���p�c���	Aq�͜�������N*�d��N@�B�d�uZ�2%���^N`��T��i$r7���
`�����-�Q6��7p�^��ލV5~�8����7<嗝b�u�s9��3������/2 <ѳ5��q�m�D�r�qQ����Qg���˸g2���m.��Ã	X�����7����O ZX�.�J�_t��TR�\!�RA��Z�"���J����,���.{���"/t|�k%�s�Cõ�U��X��s�rSl�Y
Ԛ91 va��U:���a �m׿^_���MŏTh?����%Z������t�ئBCSVA��;�*<aϤ��T��R�,!�= �a�y�Ws/���ƪ�����������΁7�ʅھN+�=���ARae���D�k$d^���G���*��h`1�~Y�a��w��7�Kh�&�r���U{���ӽ�WaSx�݁:/���s�k�$�e4;r��%�УZ�fJ3#EqL;�"��O_�9�8��&Dj1��d�f
�3�C1)f�>^9-_�R`��W�6�<�#g+t�8pm�C㺼R��j6���u�_�<$i� 8����b�ʷu-C��\th6&�{��q�˱����c����RK�it�V���ԁ�[��d���ŀ�^*VeQT�{�Sd��CJGl�A��u{���}�\�x�ϝ���L��.;?��=��q�,Rw��-Z��Y�>�_4�n�@�DFp�>v�9�Z�fW�M��:�5�󯱮�gn��l�&�h��)���l���NP���{��DK�4��;bi#&i�j�2�$�v��+�e��kB��.XR���t�ua�#��|������X`7���Z31�a��?浿�,�6t�s�a�ǡ�v����M{�Y|S���}\�*��J%֜�r���f
,�� ���[�H�������ə�,"�S)�{�g'-�#��6adO��߈V�ƙ�2��Y%"�U��е�>k�"�U��m]tl^t��/�n?LY��:R?���0p���B�0��)Y�,��p�q��a��P@J��'�!�X����JĎ_���ܿ�XYoJ,�Р�j���v�����` x�{�"&�o��z빐Yrxl�^KҘ��6"�_�<���\O�Jٜp�)Fĭn�	x��g����㳀��:���n=J�$k����Fl[��s7�`�7Zsx�eK��*��K�Xs�pJZ�Z�pN�q��U}EO/�K��R�l�JHzI�3��;N�u$;t�=^Kc ����@t��.�WH�w�����Vs��� �%���< 9�{s��gĥ��q�b[�-�Y*�T^f���ն$�w	�w���9�ؾrw�3������
D�σ�A/
�F$v+�=�=ߚ?�~�.pBq�P�͈��wU�/�9*��ajD�J� !Zq��;�k)���S�R�S,[*[�P��jP@0���W�vSq {�v�,�4���O�
�� ,y�QT\�p���pM�^�����8�Y}��=E�WjN���6d�F�l��F��_A��g�#YW�4����H:a:GW���+ő�'HaJ�� ��RR}!���.�v�5�4�YzhSc��{z3�oP��Ι�������*3��c=���0L���N���Q�o�ȶǕ��U�;���B�(
oN��<�M�?�v��u�*���ҥ�^�Amn���{��u��p�}t#/����S����	!�j���!c��_)�� �
�CH�7A��{�9�M���?�?�XP���#��$�gPĲ9_��ө8~��������!a�=g�D!:�^����[��w�!O�ة������)�HP%����Р�������g�+(K�7���������.9T1�jl�zH#�6���F�џ�]�3 Io�e�ͱj����6yS���p� �Ǎ�,�Ċ��K�X�Y!We�t��LW-��f�Q�p��w�G�72�}$Gn�hv&�,�;�I.�Z����t��= �ŷ����ʣB&ض��!���F'�ku��V4+��	N�dz7u��L��,1'9�8&�D��;��Tf�q��*?J�;b�MG��jl�t�ō��O�{J�w3�Hp-d�%'t��xrR�m%��we��������L���n�$��C���E�z��Mh<᪮zrv��r����H��#U��`*):�Z��^.I5r!2�@�$��FS�0<�� ƚ���w\�!���w!�.�l��}'߂�W)�!n(m�ѽ:�eܘ��J�A�`[�l"�Ep��1�o
P~YP�uM�>`��aN�T9z���#`a�eT����Y��H���C��h�Q�xgZ��!!B���p�m;����t�.�ҧ�.�kQ�iQ�i�9���i<�RT|�eE���}qZU=����I�Z2H�fp w8�P9�`���;l���T:�6^ �vw��P�>�cB�)�|�ph��ZR�
�$�e0�T�Rx��4�m�7�H]=���&<��5��э^�<~�)�/_,��#�@WLw��w뵤]� c���	m#���0=���j��<���)5M4��40� ce��Ot#�3��RCD���P(^���s4y �6CʗYB���&�|���fg�n�<ԡ@�#R���Ĥ��*Qt~�^�p"�n�?R��
��� @VZ�ӦDC�{�``a�!ĸ����ɻQ+�T8i�h9��>�k��H�-n߲�H���;���ߣ��0@D ��8��fߦ�@����tR�lx�P���4#[�HA��$ء�f	�2Ϋ��;d�=Ox�2������J�����!����`\�n��Tl�vxZYFL���T�@ܾ�U�&��W�%o{�5@W�ɘP�sU�ߗ>�l3qiIg��򟣿��b� �)D�4P� X�6X�"(+����Y��ܛ!���@]��m�]�Z=��ý�i�k�s'�C��'
C�G�4
��� �ĵ�>��w�bs�<H�5;��&�]8k$P-�X6�^9L��#x�G�L�Q���
�4�d�¨`�����"���>�������H�zqA��V��}�����١B�g�cŮ�㔰���a���������:n����A��#��J�@����m�=<G��Df{p�^ԟ�7��"�9\�������9QB� �����;�����!��F����I���?���~��E�zC���#k����ޓ����2����O+˨��s�J���U҅�����!�ts��2�0h� �$�
���VA�u�����S�H� RY�f�c���Z2D� �?MD�>S�Qf�٬���%��%�u����}Ѿy�y����&}���}�nV��p@�),0�� /풌L�H~1l67�o�\_I�s��k�\���Q�H�=.ĖB�6VR�58��]�X���!���K��l~2}	�.}�%=?�N��� �x���RD}�j�u���^V�HAԠ�T���-�X=�S
��5�Z�K��7!i~f��r�_~X;x������s �`<�� t'�N�;���b�Y����|�RԺ�
��m�4�p��XxO(��.).��	���%B��d�d!)��3md�(}���K��qw�a������G��%�M@Q���F������M�@�6�����r��t�`֧�r�^�4� ��������k0�z�n������ˬ�1��q�q�%0ީȼ%�G3����c�'�v4Rٯ�?w;*�@�W�z���/�@�Lx���'�\�����1�����u[3�H�����<��۳��M�q*}�RS����4 �%�`�ţ�蘕�P5�F�P�n#�l��pP�K��b��$,������^LH�O�C���� 	R&�"|v�������t�.d�'Z9i�	Ar��@���ҕ�
��J�X�(���DA�]��j"n]^ ��;:�_��%�42�� 攮oV$���*c������O����2{1��C�Y����P�f[�y�뮳y哟F_�yh�TB*o#�J�>o<w���7z>��&n���;��r��0�{3f�k�$�*?�>_�x'�?Q\[u�;���G�0QL�ض�)o+m�����@09͙G��W��;�����Bä"g�b|*�*�S�1q+~g$ �����`D�0|�vx�x Z+�:zq������Ε B�VU�lN�+IZ����°e����h�2h@����*� �'U*�tpae�p0�W ����4�
���5���Q��G6O�b�k����GX���+����D�zIv��d�|T�LZ_a�
����;�P�d�D�����~��Wr�)p���2�t��Wm�.�V"����֣F�P80}86rjJ�ִ�����9�
�t���S�?T�x��8��R������u�I�ܿ��9�ƍ؏`�Xp����>'1��rU��Ŀ�F�Z8��S �|�,5�RW�5=�{�����ݧ�����1��[�
�fbMl� N���N���Fu�%zMq?�Aфv�����f�T-
״��z���P��	��86��`��nHb�׸�ָ\u��n�\������,���S)��~�a΋�a�\��~�`��LB���3|ώY��0��c\-���;����ыv��8���/#� �
�XD�k���ų�?\��"*�X���GL�F匬`b�ߎ���1�ϗX��:R����S�|2�8��,�ه���Qo|���|S��{��ߦ�j9AmI{m��>�>�d��%�3K�
�<�"�l�z�_q5�bmyG ��Y���Ŭ#�I�'��Q�R�p(%Z{����Jz���C���T�S?�
��Rt����~nk�>�m��(Y4�
c7 �Hf�'PC{,�3(�c"�r{�xs���d9f�c��2�Ӣn&wm&�� 0�+����8��(َǨ���^�\z�~���Ҙ��Mn"B#¾/��m�V.7
��ܶ#ˊx�%�a�實��?)�Q%��*x��}��?i�kh�BU�ށ�d ����2�?�/^�n��q؃&��V��%0u�Oş���~�-k���Ț� �#%���V�U���F�
��y.����*�}3���Z}O^xhj����xEl�u�vR78!��	>�4��7�9v��6ϵ�A��Z����҆�Q�2P<���a�^QsЂ,^4ަ��+��6Jv
�.ǧ�w��r�<�d=���ma0@� ��«�Xa�K�~�Wߍd�<M����~?�膰����L�ځ��G��'L�qi-4r�E����E��U�� /f�A�
/��S�_���;A�@�1{*���0��>z2�\�WS��r�o
2�H�c�v�ɑ�`(���?�,�<�%�>���
|�'�B���������Z�R�Ly�!el=�6� ����p�B�d��>!��T!�����v�l��q��2�˺E_�e�C�ړ��i�YO0��Iq��D����#p�1�n�FS�/kh���eɕ�-���s�b�Q7w� �%~�;dp��#b WD-�	�����$�6���ҷB�k(5q�4 ��g�7Ŋ��IG�eL5�^�<�rb�R��������̙T�^�S��U��"�C�S�x��e"_,���Y�L��9�E�I��4���"~�^�xd��j�!�(5�F�ײ0�+�?W�h[$�8`,�߄]e�9|pAD*4�EѮa�Z�F�؄��q.���j�A�"W$��6C ��i���C��b��T�@��~"��c�rΞ<>�3�xd=��Y i��N�U�9��6����K�y92h��4�b+U�4.
s���D:	iI���(��Y�|Nb߯�17��}��F|��a�i������QZ T�)2����G	���9���]~7RTR��@|�1ִ��WJ�����I*��"ـ�V0�
���
�ph&_,�4n���G6@�#�;܈�v.FuQ�X
��M���6/�Xo�un8p�}����c"���ˎ��l#jY���e�
��J!�N���E�#�7a�6�'�S����&�X��}�*��J��l�/��OD��8M�� ������}������S$�ݹ�*�S� ��:S�d�t�*ƋL������,tM�R�@	����X���������Y�\F�!�}�T�n�o,g�"�o��0.��cVb�+#6�l[�N��0R0}2�e��ĶB�U�]v~�*3+� 7��b�޵4����_����B䭑�I����x<߸͆�x� ��H��H2�� ����7:�d�q��@�)���P:�j�":�c<�Z���xS�`��}n�6e�	nn*��1W��C)+�0�}�X'9������YIN
3e|���m����j @	���7Ͽ��4Y�r$�O��s��p��b��,rL���S��"�\(xq�$v�0ƾV�h=�"�ma_�CG���������X-�����eYQ�V����.��K�Y�` �/1����tQ����*�/��D���0��
ެ)���p� �%�+."�?,���������(� ���#�)H�twwwI��t�tw�Hw3�1t~�Z�O֚��g���;;����y�$| �4��R�v��������t��RBb� �lv�O����Bygu��c=J���̪$���a�2��Ύך�榞$b�F,��l@���H�5j��^F�����H�X7.�����'��'�3�L�b���F�_m��ss���H蓡�ZW�?c]�Q���?�	&]w�k�8ކUj��%~Wq��m�$e�bxKI�o>� %��O�_~��9��m,��6�����1d
n����́��Th�9^V	#3�ꎎ?�=���r�4-pc��E��]C���(�������}��E��wo'�~K���x���,�|m��ts|˘�NF[���ol���S�uw�4F�����]Ђ�0hΙ?�'�%��_�6f�_vS~I��_�*x׉��uBf)�l7��l��1��ޟK����g2���,�GP+n �Z~E��k��{/k4�w��6}W���i ٿ)@���{�B��ݵ�?`�h�S}���θޤ��AZ�A�z��T�x�͙��!�N�����qwJ�� ����i>3��wOg����j��3��s�B��Zj����#��:<����+8@t���jr�Dw����*w\�,��w�T�*�L��A�_���*��Q��� ��Jt����\y��oPX�G֊�)q��X~�_p}������k�ʺ�%:���F��t�5��@������ƒԋ��;w�'��J5�uOױ'���IԘ�3{�vP���q�5��E��Ӊ�a����.�A{��	#��^��H>;�N����6^>��wlA?��`�-���6C �ޥ)�c=��ƜS�S0#a�]~�k'�.��I<7ox�qs�����)5q���H�� >�yF+��hi�:C>d/����!��!�w4ݫ,�7��(�m�gdA�u�.��+� n�E^L��m�L���/�9:C\H���W���72s��� �)��z�Al��O�O��˂��)mzQq������I1�)8OsH�g�m��ʟ��u���A�{*k1��x=�����3ڛv��*;��]�PZ+Z8뫣Y�}�r�#2i��Ui~u&E�	�σ?[>V���M|B����ue��!n��V/z!<M9�M����l��>��v�]�3����^���F'��'c��:D�_�=��:o��5(��7�Ynb�ē�� �wj�W�o� �"�+3����68w�p֤2��C��)���{��'�x�Nc��̄)���}�CJɲ�9$<<���H"a��[�.�|	M�}����.D,��g�h�	�FZ��.�w8S�^P�ɺ�$y{��uP~Z�곗���z�{��2����D>K\����mFkD���+{?Ȏ{mO��t3���Ϭ@}vT��%`���u�{+kz���p/fCA$��Ϋ�0���;�_�V�]�)���#�Z�����[]7�v.�%V�pjn/6�0����Q���飼m�lN��/���;>~�3�����X��̮����b�����g�5���֚�{{l���Cx=�+�2X�r�v۠�����5*}�;�q1����=��	ݺ���
Gi�p���������~ty��tG���=�+� Oݜ����k0�(��=��{3�/�{P�z߆�)̆mhf�?����qf�u�hP8�s���cvĽ������3�����v�9�����\����O��������wϣ�b���Ы���r"Ȟ��:fUܻ28Ck�n�׽iG��rh#�Mi ��<T��,�{�AӬ��\�X�.S��Pm�A_x�wbx�}�����X��N����c)�>u��m��&�MM�(��I��u�ՍQ���H��~�}(�������i��^I��T �.��o&\��زRz9r�(0|ގ褧�1[B�XbM2j�l`��_uB*����lC�oO`��F�m���}2�_���PI\��*	52�枩���
i�l,B��~�@)�Ⱥ�@7���6;]s�J�,��T`�}���>�҆^��4VD\,�Qb+.�JMM�'������nC�~�w��x�҄�̂O
9,�XK���(����l��!�o�Z���6�����ȄA� ��\��o�oy��Ղ ������?|�@hU`C<�YC����&�V)I�E�C����&�1�XT��N�3�[��14:i�W��f����@UN�tz��E���
H0���7���'�t-t{H�F[Z�U��G+T$���y��(��?/=��P�8�C?K�.�(V��GX(y���v�YE����U���'�6�˲rt|=d7|��X"�L���B9X��i�H�:M�@���:���.���>��I+71`��R�'�F�U����I�[Zԃ8�
4F `��o��I�]� ��|qq��u�C�U-��=enAz�:c'�+��vY���\X�w�����ll�u�Bͅ|��S��e����>n)�N�+l:��*����￪h��Z��<a��j�����5�˪�Je��v������WPk�ÐWCTm?�t!~���/�?�1<O��2�P'B.ǎ�`����4ʻ0XLI���3�L��r^K�T�c��k&�"5^��P!m~�O��I�l��Y��Ym���t�&�Һ�I?F8X���c�����"�2�.ۼ�SՋ��e�aiiI���_]�=)�������l��R,�*��p�'T�:�����&��|䏅x)��O��ۭ�e\_4�w_��4NIi�]�����s�ōڅ|�/ݓY��[�=A`�?�Voҧ�C�ŎI|um��.�������RY�Y��m�F~)�0S12��P3�l|�"|�u�Cc��A6l�@m6\,+M��;�p�r��p�I��H��Λ�l���ɘ��+�$��q��R�L��?|/L�iD�D�vt��\�'����ol9:{�/��7�%�����}�%R1Ǐ<� 
5�C�V3P���2=�+a_�N��M���4�:a���n�P�8��'�c3����ر���C|��[�D-C-��4'8�ty�\��6}U5��X)D�I��_��7[��"��6݀j �#w��)R]��/�ķ����L����Lv�s��לk��sK�<��D9�c�����r��D��E�r�_��QZ����(���Ùp${���7�T��5�7К�}�'�x�����t��Ӊ����Vڪ1�.�@@�Ns'�E�礧�@'p�ٌFЖ�Et�	c���z:�G�)j��>�zxx�m2�~͜aB�g���ׇL=�(��0��P�o�u�[�8�~�Ե�/g�Ϸ$��� EK��7�zS�0���Hk�cJK�}�l��G+��� Ǐ���`���6�=�4��1ó�/��c�ɭ���O��}�N�' ��4blܐ�²뷱��R��"�"H��-פ �$e=-���+k�ӗ���Q:��A��jK;��j���N����6����}�9�Ӣ���/0ZgñLE����u�^�ƣ���,y"%t���n����h�6�g4	�4Q^y���'X�
WK�Q���'bVc#���_�G�5[�+%ô��0v-`�ف��H��Y�q�	�X�>���u<W�՗s�,=�����<~2�G���?�+����*�"������X�d���~/:dx~�d��-�����������fX��y���]�p;��UTI��Û�OX���e%�V�x�ԶX�<7�G�~�ͫ� j�%�B�N����4�c;uo��Q���o�;v�������5��Ǘ��Za;Ul�jd��"ە�7XL�[�������l��ٔ�l��]���ژ��A�i�m�2_n�4&��y�qy�����g�PߚT�02�U���}Pџ����+������X,�e'�N��g�U�Y@��&+S��lw~�V������I&�'ҏR�C��.���ݴ�A��Ѻ�"j�f�]Uo����랿o��.�o{������9 �^T����Dĸ�P�,�]Z���r�?�!,a�W�yS����J���V�J�������s�>�L$_n�fm�$�J����S�ݥ��5k"�Kt�uq�zqt�*` *7m37I�6G��9�Z
�wH1- ��� ��ES{�*������t~x��-NҮ��G�Иu'�\�-��/� �Ob2�w�SM��7a�P���,#w���+G��f���]ל�@D�틀ye��	�X�r�~NKSReo�\CE�Q�V��������w�]�jq$p��.N�k��v'�s�աoك-tt�iM?&�rl� ;��	�-�Pz���*�n��?�* DmG�n�+B}Τ���ar��F*�ѿ��_>P�f|�Z�SQ,:��1�L�[�7.J��U;��,R({�S�{U��y���d\a|��g���'LP�L��}r��W`E���\���o�����ܚ�I��.ٴ sa�y�g���rrdC�Pj�:����]鱗V���)G�P���A��i���9���v�Z��<���^�=���7�$���:s!Qg�n�� w�����Iq�N��m�*.�n�r��͆�)����{�/�OI���ZT���坡F���E���o��K�.�F�duGM|>|i�)�Q��7�����w��y$�~�o'|������Л��d'+EZ5�d��^7��U���!�����@���G�����\���baڊ(R��N�>�<���@����b1�
޸���а/ �w�V񭪴RD&� q�|;�-�=y�z�L��'���,�����7f�SzS��?��(�I��wn�Vx�F���?�C�O�j�i$%��W��Ν���� ���qcv�D�TeD�?�%���yʌ�V=Ln�n+�WMnQ+T��V�۪���j�")�f1d�9?��JO��<B;()�Nގg��C|;���&oAtN����n�s��ګ�Zr�M2��xo�§�����Ү����BC	AF�N+�+5'wwKyC$�f�MJG������XK�"�*&<��[��d�_���9��i���74�Am�;��rf���13́u���n���\YR�V�y��l�F�qr�`�ң�Չ�T�Ի�H�i��{���E�z��V��YU������"��~�"��DJj
~��2?Y6�"���(9�g�(�V����:��Ұ����1T���Ԩ�_���f���\4�� �2�g`q)w\%��5�S<��:�g����m�[����O"�G5�J��䲸�)�/<S'����J�]����KIS���[+�4�Q}.�gn=�
W�:�dҪʉ���D�ț�M:޷ H#F����d!�����}ܸ���>��`�d 1Cݭ/7��y~rE���fx�������w�)S��ez
�����z�����Ao��=��+��+��p�~���6�_D~Lx?}�fs1�? \�IO������H�8�sK�E!68b?��Li���𼌀-�G�b��BGX��t�Q-ĵ���������Jf� ��;�����>V���wK�X0C����TH�M*A�|�S]���cļ��?̆�l�\UI$��7Yi��e�>2����X�P<r�B�h�,���2F5n��0�0TT��UJ���w��
]�퇙E]���S��5�ld��_Jw���|p^5�)_��H��WC�'�hѷ|8���%|ѹd�>p&ӵ�����跈&1�$R(�5(��@�QH�jq��fٖ\vvD�h9��p!`�/��k��cX8a���5�-�.��H��Dt��=�/w��HT�[��8��@&)�oq}���u�W�y
�8�={��aӵ�{��lU�E�C@�m���/8��67�̶t����a/����bqJ�t��bP���{��%F��P�~��2����s|�n�>w'�~��F۷*q�c5Z�>��8.�'P�v/�y�
wT�,�N_d�g��0���&N.X�y����(H�	Z;ÿ\`���S<�E�n��z 4�i�'����Նwӈr�Z.Z̉��4�|����I�\I��C�u7��Y��CW�@-.םr��3��ٽ��m��y�]󒱨�.���t���
��ٚ�#Sie&�������c������ht��3R����r9�>�D�~r�J;��'���B�G�	;)	:�G�\m�.�d�����lW;X�3�o�о�(�"\ D+!���:���bZ��a�"\!__eS���8����0�A��{K�s�o�?ݎ[�X-Ӧ��bCt.@��O�U�qi̐Ά�LO�|v��g�w��/9�C��Wy7�u�*|(߱�e|K<MrQ��e��b��2wآ���yA�MZW�g�������;� ��,�P�Su��}s�ꪚAE���U�@@��{^s��S��
���0�
xX"�3�Pz{*�Wy��~���7�H���e��*�����lY@Q�]�%]��rN9A��m��2��o΄hW�5��1^r�>��#9#�'H��&���}�լ�UsB9L$\�1�5��n�g�\`a�J"2�n�o�&ZF�Z�p����tB.y��>�ݐ��@�����z,G%���0/ �P[KLӶ�H��R�CV�����e6f�q
m�Z��~�tpH[:�lf�!/�0	��� �x��a�<y��l$v��= KA1U�U;���"vi�nU��܊��0U'%��!y�q�C�j^,�B�T_KW���\76�o�F
�0v�H��O�ԗ���j���
JGl�˟�N;����PB���"��D��8o]6�
�ް#�)�l_����P��s�v�sh�1@�ٓ��.b:���Na�d�
����oxd&�eSُE�%*��n�+]K�H��I;5nW�(������ۖ0��h������&?�iH��u�Yp���,#��\n�L���� ��|=��Sdm���>ͮ0y"�@��K&�V�����'�W/<�����&�/��z�?�wg����F}�Ņh��N�_C��j�Ϳ7O�#��&��G+�q$B&[Ԣw�]7U>�=?��.?w��b����B�q����'�������,��ti�"���U�_z��
�¤�T>�@ϛ�}Z�.Wѿm��L�s
,&d���K���L�E��zհ���~詍�����@�^�Bl�ۇ��d�Z����/�è.�,9���Ade�©�e�(svo����P6a������ �F�@�����1W��"l��B��%/
�
���܁lO�Z�>h�$�Uy�h��-(�`M�m�sQ�}\����T	��,K�%Fg�R��]W����ƔM�+�6��v��y"����Ҹ�,T��u��tb���G&��}�HR���Rᶉ���Ȇ��G7���z�"Ϣ�
���7<4H�jz�y���A��߅k�9���}7�=Ts���v�+W���n��~m#��&�\k�L��-/�
���HQ�6`a���p�I<DNɈ(�hJ!��m�!��G�	[Q���_ku2g��@�e�T;����掬$L�Cc��b�԰�ޘ��P���q)3���h<v�U���D�dt��3�81<�i�'V:��,蝟�
�ǎ�����=f�/i���x�O��
��+by�=���U"ߦ�ު+�a�|	��=���fG�ܢ˫:A��7��WHx?����G���t�-iu~�%�:��3��6�#p�k���v�bl���xa��;{��Mݛf��@O�zT��u�O�Ñ!����B�(@ g6�˱�dzm��i����Ո��_���3{��[�0D��暥g��fn�#!s��n���&��.M�Lnl��6K���n"00ߎ�jx9�4�S9�RW9;���y����F��?w�7*F�E6�`��
d�5������K���q؛1P���;�V��K&��LD�|v?��e��4ɼ��_ht��%H�����fG��e�[TG�L��xݜBlEo���xd���	w�~�Z��/�����_�'E��^m�t�i�qx�	�����V��4}Ow�".>�B*���N����w�~w-I�_��e_�4�������im�%Y�!楠�?�����2�}�4��+��i\�ue&��,5�0T*)v(:�N�d�]��=�q�j�<$�@@Ⳉ�T�ÒC�ć(��.�|�R0 '����>��;��p	
(&��9�}�G�\ 9�D'�zWm6d͙���:��D��Ԣ�����3�"d��7���b�r3=6�������[4)��� �v�Kg����v��4�TJ�O�c�M�G�<b+��Ȅѕ��ǒ�qxZL^sO����vj/���I�aߦ�V�+���~^����B&+.�Q�dV�KݏY���j>��j��(y(4u{��Ut�4��a6[�N/�i��.ǲ���]�~sq�&��8(�΁4�me̗�&�6|�ۅ��~�����ϼ�BDW�ӧ��)�|��G�0���	��=pEiѳ�K�_�V�Sؑ��z��MV�.+�
fym,?[�k6�(��ܤç�㯮�&��6|./�T׼J��9Yt]to�R���mpR���{I��L�+J"�y9R�h���i���Q��l���#�L�9�Q��:��s��"�У�m�Q~f�	C8Q�����\�yC-*w���߭M��~Ԋ�����x���m��|�`t��3q�5u��U��j�u�¤��x����w�y^�x������}" �1��+5"�Q̿J�I�L�Eu�)b��\��p^��-�X��pkyp�Ov�-+϶Ȫ1��EӐd�y�Q�IwQy?[��'��	�,�Q�o��z�/v�_l���*�#o��g�v�����b�u��?rp3 g��F���QMS~�*FF�W�W�|v3|�\�&W`��TB-?y��v�uՍ����V�=,��[}�9�֨��I.�t>��2}׊{Ӛ�E� ���r�B�S3@T|��| �Ns�(R(_X`�z/V� ?( ᳴�o>ӈ���,��n��c�,y���+��O�������PZ�tG���o�`�೓�/�j�fzN��� ��<�]j2��vw�?�n �1�h��4���.��U�h�|ƚ�
/xѣ���a�
Q#Ã�'���__�>8��4��w��*�n��R,�:��/��%�]���5jJ k����v�Ř�[)D���Mb�:��է�4���S���wK� A�2C�ᙠ�j�a��w�I �\��a�@�ܡ����``j�S�����Ƚ^�?���V��yl��]>v����7��{�g�1�bH�aP�O�n�%0\��=�u�}���A�og= [���3��b��;�sr�דJ�YA*k;LY�R O4�a���dX>A���U6�3�V~���Y=��*�i����[���^��y���A���DV�rm^/3���afyt�P�w>��4�dR�F��=�	f�	j?5�a��O\�F%eh�ro�sH�욥uիʭ�tXgn�g<8	W�G\2WU�*a:�w6�B�Ŷ��vB�1ĩ��V^�.�u"�������|�ղ?���QKy�!��'ˁ��f�p<6�a������K<����d$Ý_����������x�P��gyX3k��?bC04��.>����9ڙ陽�}8�<N�L�ɩqL6�~����n(Aԇ�(@׮T�-P��n��}���w�=�hW��jPC�,���Chl)@�'�vU��;(_-`�dW��S\�����tc�=\%�I|f� >z�"��xۇ�wvD�?C��4:�m��>6�ߺ��r4O���U��[���kg��p-Hzj;�GTFz���^G,��x^}�Xڼ��z$Z��4"A����n��8��-���j1��5�X}�sk���wg�l�;~_���Kw�]����H��տ5(�8$�}`<͚Q>{�} �9�Í�~P�aTb����"�������B��s��d�0�R�s�:O���������y�Ւ����~6�w�aP��A3g���o5z�=w�L_�it�A��t�I����X�T��f��~���}+ ��X�f���Vk���|�J<d N���Z�F=�-��pk�p�;v(P�^m%l�E״���{{�S;4�<�^j���8o{eü��P���j������@<B^+g�f�k��!T�O*�$3~�kڲ�=k�=C�"\ŋ��!4�v�s�����f�fQo�~x�yVq��d{�V+��;������/?xc�Cŝ8w��n]fpkX��S��&�*����z5��>2��ۿ���0.�w�5n�����6X������������}�n'U����<�b�|��#�X�O�K���<�OʿW��S�1�
:}I;B�Js�K)4�:v��K	��x>���.��nh�����b�!�Nˡ�J*M*��'1�P��&�Qw�W[�d�J\��ʻ�R
�=C�DXF��e���B'	�s��
?��P�0�Ĕ��?�����xd��є���+�$k N�K�A�zT�N�wp�bio���*kl*�Y��op=v;��适�V|�bg�k@��Po��@�� l�����w��>�	9Y��|��S�6;ҜH]G�k��y�S�+ٝ泍s�
�8XKe>���n�����$K�k�g�Sc���&�aۺ��X��.�:��}fs0n�Kw>���l�(zd{��"\�H�ޘ�ӎ���uyT��*{{�K)y���蓈*�N��\U�-o��-^�8O�pbc�w��3���K��Y��}�u�Y�NQ��f�lv�=���7��5SJ�Ka�ru�v�7�t=��`��O1w��ZP��-+ I��q3�H�5��g�Dt��d��~�b�P���/q-"�E���9	ݙ"+VD�B��)t�P.��邿���&�Vb�Gu����e`���_e%8��L�=�x��ax_�T��� mJ�$�����v��gC�������������� �����j�Ϋ���W�#���O�"��0���X+{9*'������n�I%
�Nv��H�}���+5�)*�>����fgw����ٗ�OQ�QlzB���`� ����_uV��U-����; �j��"�D���p7���@>��>��^�~u�)(y	*����EĵC!�Ӷ߿�1��cG��^#�W����hɺ�亣20�l��bg�I��C�TVX���x��^�O�gJx�������γ@!:� ʀx�Lau��!����.=ʕ=@@�~�s��{������lW�	/t�lO{w��2bE�wa&�ђ�!V�ݹ�����:	`a���p�Ĳ�=�qI�CJϴ !���0��i��I��q#�qf���qƪ�5d9��ҧvŌ��!��N����P q�o�~�D��I�LО��{�M2�������/CK�̝њO�ǘ�\"�/ RtB%f�l�h�(0��M���;J�َD���F�ˑ0�����+*�%ĵ'�.���q �V� ����u�rv�X1�b�J~�oZ��$�挎:���� �r[�7�=�����C��*f\r���R�A&��^}:o#b����r�Yk%�y���:�X�l���5xxx�(���!] ����n�^�vL�|�iLڍ���'m��8);P	�a�����!r�4Ek!d>��V��4�l4:���s|��� ���Cw	�>�5�%[�%�����q�X'e~�����I�E+�+���}���7m�VRX��_s��X驙8��ͫhv���b%��9S
���vt���撷ݿ���X7�&�9J7i^�a4� :^�I(�䇟��N�%8��G檄�eИE�zX�� |�� i����%�Hulf�H�X��o����5p]\�l����q	g�x�+\�Y2�#��c�UЛ��_xP��
�;�#L�P�@��pL�Ƣ��i�X�k�q3Y��9C!	ty+�_��G5tޢ����*���7:("��������3RźY$�o[t燀Dx�ߧ�LH�>�r�ӭ,<ٞ���:�mI�1]@�B����Z�G]�hA��|x����B������_�"��݆"�B<�O>�>W"\�w�����ie�_&�f�ݭ�y��M҆��'�~Hc	f��~�v�+,��8��n�\�=�C����"�-7��.V,���TG����o�0�������z��c%�3i�>�����Izִ	���VҰ�����y+?���nx��	��2�w�?�H�Е][���4��1�Fg�>�+�ٻ�/G_ �x�8��~�T[�4Bő
)Ep�=V��Ŕ0N���g8�O���1fl,�>�`��4��bw�߳J�jXp��E��U�H�iRceHB��q��n�F]���1fPm�1����� F�"�w��}ֹ̮�����R;@��x8���K._�E�7�������U�M���+,�$�Ǝ�j��K���"��:��Ke�>��W0�x{'1[�����I%�KM%I�a�)ҵC�!����훥�L�8R�*�_�D�JIM���Bz� V� |�$��agѺ�v=~���yX鮌�������"O�]��}���I��<��0���W�H�䃻8z��ڞ�S7G���#D�졡��t�5U|��s�1e������t��G��f,x�l��׎Y�7�#w�+m�%]��aL���u����������2��n[vt��MX�͘�@!cH6�<����wkq�>��xo�W#vQA�",����6 j梘��X���vCd���	c-O��ˋ��+�I�zJ� � ���^�&����&�y�����
�+1���O���F1{�z���t\�K�/�V��
x+*|�x�t$��mk���G��	ģ#1O�����2�
�%��[�i2X IO������rĀ�E��_�j�wKa��:���w)��+�~�V����&Q5�q�)͟N�K������hy���f ��טq��LjS_�����?l�L��݄��	�ލ����Wo	B��c� �;��o9z��Aݨ|�c�
<)����q��`��0��D�|�ԙDsc<�jX�骂\mC��B��Iު���n�J�%��Ո�#�y�".O����jW��+�a�t"Xd�"i��T�ـp��P��/-��}��N��~�XB�2DC��Yɚj��L]I�v[9f��Z�Ԭ��^���)����&[Hd�d�]�G�r��_�]���.@q�$\�a���C�nH��O���V@CK���~��	��M7���|�o{rp�]	|h"�� �Yz�,@U�$!���Up�Aw ��S����$�KO(�h�����Iolr�c�<���L	����'h�g�����:�C��)��fu�ӈ������e��j߃t�pj+}�5Z-�%H��zU�R5�L*,ӡ*wζ�I�J�b>��r�yan4��KX��#;�Ǟ�Pr\�7V�,n��"���2F�h�r�w�{ER}��q\��Ws4�OF|��:�pU%q��&s�|�\��4ks�k?� ����~p��ǆ�]��5��ey��JT2hq�c���	���q�G��d�/yo]Ȁ�sS����������)�%����=48a�v�.L��«��,sc��#W��`��Ӂu�!���0��_f�<�}�u�n���0plgl�uq�B+�I�(�qbK}�K"��g1��Q� �Qf1*�Kn(�:�ٳ����)m��	���I1�����@х���L��{��7�~���u����xAn���U���3�K�A���ս>�3����6� ��cf�ݏ��Qx"�X&�y�z.qw`l4|�+m�l��z�z�z�4E�pw���ng�ux���#H#�pF�j�$pP�3�;�Hr��y�/�e,����'ː�'�Y�`i���_�����\ۧ����|���Ř��;d>W������\�ԾϢ"�>���t5��߲�p|��)����d�p��͜�X��ou<����:�a��}s���6hQ����d��%;?%��ZfZ��'N�asni��B!�{��|&8�����yW���e��4Z�2�ӷF�H,x���r�Jr>W}o@�� i�eU�}�H�*�(�$jE8�|���z.4Y����@[�|�]���FZX�ls��P҉�=�tq�~��:�a4�U�˄�T�'��,j���U%�|F��S�|{���;����]k�Yy����ͤ1��oF�r��~����`������Zl��q��ҧ��/���w���Dh9�^\����3�)͊�R�E�f�;��\�*E3�ƻ������E���j�N�,�ՠ����U��)��=�hqa_�q��ϝ��]���du�[RՍ�ƌ�ZPe�fpM9K�S�e|%�l;���q8�.��L���S�OvQ�,O�Rg֋�s4���{Ai�(��o=��w��	C��t.F��ws��b��&b����.bޕ���ͷ�	��ZF�3S6��	`���s��S��r�RZF�/�f���Ț.�vP��Q K%&K�:�&PZ��s�)��_Lg[ZԬ�O��9�^��I��u <��$��H*}�U�~�A����/�?�=T���2��+�/vWJN,z[�ǲ,K�k5ӹK`�a���
(�U,��~�Z2V�/z�53��|��%�����I*��Ԥ�|oD���Ru-���1��O6���n��QLZS���>�{�O�������VL�c�����x^�r���3R=ӸR�.�x_�W�b�o�-F�
�YxT=Z�ʱ����rz[�T��sdׅk�>�n���"�iZ}*ͽ���G�����2&�y��7F��م��U�B�附�J0h��XW)��֢3���S�2����J�&�H��WQ>�j�KHo=g�:��e�<��'���n^}�y�8@��:k��]���bi��0�\ٗ��s,٥�cx��3�W>�+�i�DV��>���8�2Q�p��+������eEK5�*��םc?oy�%�(�l�b��(9�*E[K��E���B�>�w���fm�>> o�>���)�Y�ˌ�&���U\�rK���ʼ����c5�V�H�s=�N���������y�b����8�˲ٵ�w��Ŵ�#S�{�5��*�`B��'IJ5� ��X %��q�V��{ky�n�[�I���\\Jb�`P���埍�D=-�^��Ā��*��z���Y Zѽ��T���C]n�Y%�d\�)1%X��3��,������,q�_�A����_�zrwN�.9��	h��v ��1������z�?p�PǍ���2�w�o�Q��#�_-1ȌE��EN��{��ݨ'4.֋���[D�0�&���\��I�at�Wx
�iI7D�%��X;=��ɸ?�ؓa�K��l������σ�+�u�O��z��d�
�.�$��.�g�1ث.6����z�V,Ġ�V��*=�#�  �O.���q�ȿ�������W��U��}��O�pE��l�~qF�Q�b6W��D v??^��g�#�_�Yz�4LĦb�� �Mj��`͆��평@@�*,��Y������,�䷖����	#Ũ���Zby2��.'�!�Ӽ���ӛ7!'���&��0�F_��v���6qP��9�c����S	N��8c��E��T�4�L���8A/R�OB���}��o�0��U����<�F(�<�#�0}l�F�=|�0�����MyQ P�Nu ���η�C*U�N.`%�욟ۉyw �-i��[7�8q*uC�����)=��&�� E��H�J���fZ]O�B�0{a��U��[مl�!~�9�;�Hۡ���Y<c�m�k�0o��G�f�ӫ��?�6w k���2���@b�5Q��JL2���!蟿�[#(�QZ��q��HЩo�ׇ0kj��:����_�Xy�9�w+`	�Rf24����GX��e+X�Ɖ���~ ���(Dqp�~X�ʇ"2X�|�%E�Pً��Z�i�X�2�ްrXlo�y�5�N����>�A��|
fe(�#�o��=xew�P�i�AU�$R�_����//�Z��f�\M帑�nsK3q}�Q��yW�"�VAn!�3��e4�RG|o�-ս�T�'�yx����̳��tC���9U��]`ykh�����|� r�Yenw��{;B����
�0""��4gm�L1wt�=8����@ q^��(7rY�?��z�TZwX������Rq��	s"*� J�"B�� ���t�j$}�sWw�sJ�Z/��ͧ�DZ��*����U���񁯴� ���GF����Kfͮ)��L%��D�ka�x�zX�E>;bmn P�*���[͋�.G����{�Ū~���2m���ZT�*�/��`_�?��e�%f�0��� �����X�qZU���A�Bl�Wp�wu���V��T���%�t��[9[���Nb�WV�Y𵁅7����¦d�E�O�}m>�]�IϚ�ؠw�rUwPKӖ��e���*��|8.S}xW#!�5�L�,˼տ1�9�10I?4��N�=�7!H~��?;'soր|����%^�T~d#�kWg~�� 0��,$�?��2��e�A�[p���Cpw'��{��!�������!��]�������#=����5������j���V��UW?��]���E�ԯl�C�JJ��e�����}	����4#}�I��1b �f�c1�LNĩ�6�q)_4��Q��5Q�"���60rf��Цu��g�Q��u?�L=��~��[�ji*�Wc�9]�>[�U /��-�&B�%�X�0N���-�n���jY�k��WJ�0@囅R�U(5��]1`3@�J���b��x�Br\;�>�S��ᖈ�殽Mz�qQ�K�\�fK�=�Hn�D|ګ��� ��������]W��P���z:�jl�ɥ�i/���N
��{�MB�ۺTh�?��E��M^"j���O�w=m:9�3��x�$O�߿	s�zr��:T���ǫ�����\K�#`�W�=v'Bkn���S���Ryw��6W�$�Ϧs{��!����.�J8�= 
>��(C�kQ�����o�������n{��JO򄹝6qń�o��b�%�gv糛�52�Rn�ǟ��5�cn�fir����\�,�Į.W8=sTΛ\K�;8�S����N��~�l�m1(��­�=��W�̣�y"�����ްy��i�!���X�r:z�1�s�+��V�N���:P��}�ZX�8o��\�+�	17O�+� �y�.��ҙ�Ӛ�
)s ��)��#���t�Y�y��5����f�/H#�2���\��[�S�t�^� @�Y=�jX�F�Wfs5ٱ�3�}w��VZ�Ja�{[3M��ە��s�O��+�6o�����з$Ɨ��"����Ő@�eM���{��o���ccd���jb$v�+��6v�%T�;�����DY��f?*��\�IÑok�Kz��E���Wm�8>I�l�#S�A�m��o�Ud��ʯD��@vN��|�`�iw�]��CRL�{��׌�B��/w6�ܚ,�!.3�<vVSr��@�->v~
�	x>qz��;�DvǇt72�>�f2
��$�����tg��XAy���rOb��T	�kO�!;�� @O
�]��� ���ro9?��ML�'�^%������V�*�l������j!g�vʾ��qqg�����A�B �w��.T�%�H���~t{L�:��:��	;"+F�������Jܿ�kn����4�]�	x�l��8���E���R�@ކ�MҎ}��tޣ��%����<�yOu�����;S���*�X�6��c�Z*��Ҩ��:y��ɭ����`�9��݊>���z�-���X��L;�Y!�š�� J<z�z�V.��=�Ԧ9�Z0hK�Ӄ^��=}I*�o�R-(R*Թys�Q��"̇lS��[}��d�`/�.�����8@�٧��n��yfY�h�%�6%�H�Y)��y�7�XtƅX��㬊m��)���߯_�[p?�O)�q���W�mO�)�E�:�
��.�{��j�.
����(Գ�Ħn�'�Gb&�/v��ୢ�}�6�Ǽ�"�P�*,��$e
0�����@S���m/��l� i7{��`j�W�4(�έ��D&�2�y�ˠF����#S9��
���%�/�gbm�6!;v�y�w�	-�)e�<��~�w˯�yEГWE�J�{t�N��p��-a���i��7��֦���O�13�Z��;n_(t�7���S�WJ��������x��,p9�_E��I�dP��<��Q+�������������fj�K2MP���B�s_g]��'v�7���z���Ϻ����C	��kb��s�~�[7�˾��X�Ķ���Y�Ht�����v%&7tq~�9�������Ga���/��|�L���0��u��1�O#L�]R]�,r��h���2��H�½�)}�K��d���4.%�������Ħ�y�v��������������*6�>���=�L"im��Ҽt�@$�e�G7����������f�l���J<'�+ץP��&q���N�iF0I��;.|o���7��3��7��_ϓ��<�.V�����Զ�-�z�w�I2G��ƈ�*�3�S����XaCO�>�(��fG$H���2�	��ǝ���K�Y�����/�yy�]�j��I3n�Y�gm�K�gd J�|I�W��3�p�t�Db��Lx��i�h���_T
v�3c��ʵ�}�I5H~?�ޡ�r�P�Mm���5�*>\��>4͈�[��v��	4)�&��\����`�;����d�NUٔ஻$*g"��ϵ4����v��i�C��Ш����zA��X�s�T�ZY�������?;w
�묨pc`�g���BQi���'�w��̘Dַy���b�)��6w3�,�����om��������"	��>ȜMf%�y&��H6Tj :�JFH��]��.������nr�勁��BXm���Ε�Ґ�����+���I��<Q��`,'���: �l�����[+G�m��Z���J���I#�w,T<�����S�G�L�j��NVJ�}�k���./Io��n�9�sQ�p2��NҷsW��I�?�O�0A�s�,z}�P�Ԗ	�L�Z�b��+�l��w�(�v��oT�ϡk��Մ^wh���0]�Y��*�ZMȕ��a.��gw����˿�.�dʨ�ߠܝ���c�]�B���Ŝ�8��a3t,kh�9_=P�L��6b��I&O*�6_2Ե�kW�99�χ{��O��)#g���PJ��6A��i�Y��/�lg'�\�w����.L�>��FM��HZF��Rx�*Ŝ�wVE��'q�/8�:��Mw2���K�"(A��p��ٶ�ol�S:�_Fԝ6�	>�we�Yk���;�D"Fw���ʼ�w�%>JN!����(�;�E�6�J9�s��7>��Jg�R!Ǩ;�B�B��k֊�[���+�;D[�-;ֺ�����Es��F�s��ࡃ8C�ζ
�.y����I>H�&k��sq�֓���INR����4�U�T����t@UO-��C{f�9����uz�^�EF�xg�xkj'��}0Q�.��6G����TDM$��Kp}]<��b�ؠ4�V�b��[�Y����<p�p�y�h����I���D�K%��`���
��.^L� ��'|:�6Xq9���k/�i�+L�]�;ʑ��)��u� ���qA�kW(������y���fE��TE�Ƒ@�lI�dZ� �	�>+:3g9���Z���ҝ�r1C�\$� �wp �G�5Q�<1�X�Xp�y�k��j�K.H��^&�Ȑ'_G�"��z,C��СlSZ�^�#�X�7��E��* �d�$ǖ����"���at!(ïu�������Zl3�6\Q�f��n�}w�5��5I����F��W �fV���3=o&�r����o�!�S��jѯ;|�5���`�'�嵇/%�_N�|ښ��/�h?4z��/��8����Y�%P�P��oO�Ȋ'j0�m���F�Gl�#�	��3��<��u����V�	�$یj�X#@d���X��L�<�|^ɮAڤ8���,e�e��|!o�0��Zej�|'�0�Q����@���-E0�a���3����:�I�)N�:��J�����6 �Wsi�jP�{� Ǟ8�ksLK���J�T��0_�ꍼ�O/p"p�TG�Fn���{lY߽�׉��&ڇ��cE����hW�o�2i�IzAÂ��c�z�2S��&"��	���a��i��y�7��gm�Z=�c�g��J��h�a%�|��kbJ�� ���B;���ڃ���N{��G���5i4��7��@l&(���1��5�{rj�����q�w�bVfSp���Ks� CJ�d��]͕�Y�Q3u�9.�e����8D@͛�}�oWh!'{�u�Q�(��Vn���J�h
Pw_���`���% ��Y���3���ډg2��G���D�6��	��[9����t��
j*�/'���w��8����!�֮���ӿߠ(d��v���4|��\�\���-Lm�g�H�u����R�OꚂ:�O��2�lV�w�
���C�I�����\�#�%:ۼn��z&8��Y���upCKO��
������L:b��F���P�A�@?a�p44�j����/7@�*:�S�p4��Xt�FJzJ\d���3�`��^>;���?<���d�ֳke:��ba���c*,9�"q*��g=��$�mc>b�a�
��	��G��=J�RkR�0�xX0u��0۠�����6�����'��"�)O�ACۯ�}���+��ϺCR~zΎ���/�F���Nj��Ȁ_�ʙ1%]���|$��i���)�9O�L9��?X�1�aEau�����HB>k#ݿ�����
��g�29����s�Quڤ1&wiYTG韷�f��)���b�J�_����}��iHtY� ~��&�z�y��x"�(J�}�WI�:K�1+�R�W߉٠_>s-��?��e���Sp���`���#)�j���0�2;�h����ih+��-��"J���$�<�F!�ǽ�O��~���ӊ���0����s<�aQ�ȝ�w!������m�� W���6o�w�D
�� s���0�x'�������� �o��LV�x[̙B"�'��x���&��&�@��}����@+�0��`��'�%�f��"��~���9��������M؟a	�I�����*'���M����Jب�I�^Y6�ݪ5c���w�(�GM_W��Y1�S��顕-�f���ԮMV5�J�
M����6e} ��`��_�cR���1��ڇ�Z��}%h�A!6��Y����>A	B��R\������,4�l8�4k{N��x�?�B~�����j����q1 ��% ��LK����Ђg�B��D	�h-7��jq�Ҷ;r���G�ɹ��̪,�����a1{xͿ�ڱU�z�*�/{�"z�Lٺyη0:���C�ڈ����`�����})=��z���硴���w�+c�~ n�Ն	�r1}gu'&|v_QG.�/n�I��`��/uX+��	��]%?&�g�+)�պ���E֍��������Oi5M��
	��z�O*�OZ�i�Y�����	�t��2���͡[^vu�a}�C��z~�m�͈"��@�t���y	$?C!E�bd} ����c1p�U^�٥qk���/�k��(�~ђ"�����aS1�N�&=eE�BI�(���=2=)Xi��7w,�=(�<�Dei���&�֡�i/���˽�hFydI�Uێ�_@q�6U���3;�cG7u�+Z��E����� ��̒3�����3B'\͏�����ӕᜯ*��'�x�M�0 Z�y&+��!g)�\㊦  D>C�bL'w\ b)���@LGi~9�>�8m���q��c�%{ݶ���BCc|��, ,�E�����Mua�{\�W����^BvW�X�X^.��E�81?��9wo�#*�ޕ��ݎ�Ǝ����ҥg�39s���,!��x���h�h}��h  �����'�o���w�v�Pect�(6%	�Xq���c��)�.VTT�3$7�E���ֱƌ+��nS��¡-%[�R�$��0��8@Q�󸒡��K���_�a��ӭ���M���x�a����a2�ѳ>�������|��ʮ��:Yb�s"�uoI.����FO�q4=ȐGbax�E+� �����b/Ɔ!oY�	�n
��Kt,�o��$�7A���;'&5�E�� �f%��%?�T�}���Z�9��z�f���E�e�Z�iy*�o���ԗ���70���˓�2 c�Ou�������Y;��E�gT�S��=�+]����u�דKW��B��!\LSP�aӓ;ٷO2ν(��p� ��-9��΀u��&|f�0$d��)�y�;�����-R�pgn�~!�=�܏ �;H���g�d)�q�ԟ���J�c��@(�����4�ɫzj��@N��1li��"��߰�h�I��ł�)�!�'�aZ���_疪w�1��#�|p��F`x�u"�+p���~�CR</=��"x�)�t�ÏZ�M�ݨ�5���1�qµ��d��B���(Mй�Ԕ{�F�
4H �!���\���s����C�E ?"��`ˡh�2��)��tL����n�C���P��G͋O�f�x��A {;ЯP�X��g"���U{m�O�/���a�.�3(5���7�^��L�5AM���5�m��v%��G�����61�ςF���Ur��"�	�>��^T�D��>���ՏIS��h��^��eh��/G�X�+q���a�N�X��*�䡊4~��*��h�{��T�E� ��t"�|/�!"� ^1��d�q�o�)�r~w�{t��	GrM�_����
�-r�����,R����_7/�4�l��X!�g�&Z�Uv����xw����v�W�`j��N�|G7��b�G��zϸ�KT V�<��O����0gM# `'�3l��A,��R�{`;�p#~֢��S7>�n)H l��K�(�KJ�)�ϭh���N9Ϙcu�[��^W�p�����5�Mz�dKm{�m8 �T�d:':���|��dA�2���!���dt#�[S�Q��
^8T�\�M����_(b?�$ ���_%����24�ɨ�D��o�����F�Ő���h��6��S4bۺ��@}g&Nԯ"������6��/ø� F����n��o} ��6(�#�"3H8?��)��>n����� �+@��N�U/	0Z��[����e��1#L�gIYh��_��Q����9��/�E��0k���j�P�@�����Yn���]�/}
�9*}X#}=r1��S}}���ڡz07��xai�ԮV�ú����a�f��v���ZW�����!H��T��y<��4B�1���uRWl6����Ko!�S��K��9�K!�mzD�-t,T�/�A�Wn����E[w��mX����~���=��z�0)%t�[�p�Ҏ�O����|��?ߜcݹ�%��������3��Z���mJcؙ�je���J�Ԑ�Q��~���i��*|�	���&��;����ב��a�0��U�W�\�C��:��a��HK%��u��̒�:�+?�P(�_�X�{"a��3�u��(���k��n-t��_�a�6T O����i6��Bi�g	�X8F P��$��'��{;0P�����<`�4�ڟD<���hcI>`��A�W�hX���A��@t��i���^�H0Xgg>(@	�pĲ����(cw"�����O�F/z�CSǛKX���4��Ӿ���
���:B�7��	��<���E꟫\��/�0el!�aGu��7����N�E��,�<�{�5[d��K��>F���F�&�a�҈���0 ��H��M�r�k�(_�(��q�ጦ4i*��Y��<dȆ���#�B�OA��r����2�v�H��{�Y�����3�Hl��t�~z��4!��Ƃ�J�ퟎ�,�,
�k%;������l;��C���t6(��o�	�f�8%&��@���ث��y��o:\��$�܊z�"�y���[��zd�X��&>	��(I� nL;��_����-��x�(ecq�eV���_yO%:��n.C��ɹe�O�k�U���]���DaF�?j�1���r'�+��#��+�oZ���-N���pU�۵��=6�#��!�!m�k5�٘z6��g��淵��|a���*I>n^��|!���ϰ��m�;���ml�o��R�Y�r����?��H�!��cb������iG�5��p����x��hQ~f^+��C�NA��3u�� �}s�0A��Q�1MC1B�;��Y�{�3��5�lMRݦ������o����gZk΍�ES�:l}&>��Ȟ3�����E
�"�T>��ϛ��ڷT�ջ���:ɞbbSŹ�Y�,)O:�g��6�W�
R&�W2�ak�h(�fl��
�h��D���6k]F)�X=��ʉ����V��s�Re��ڰ�i���I�շ�Mo�m8����nG��,v��h���ke�sXPr1l׬�<��� �H��i�T(��d׮S~�ő�"�S+��5fMd_�h3n#��Kg]m"%���?N�_��!��Y~�1]=�y��5��qbq{a�k����-���n0���o܅LT"��>�/�f��5�.���3��yB^��>9Я�of��B=���U���5ۙ�幮6�ڬxB{�S֮;�*�C�����0Rq��h�׺�q�qÖ����IF\|I��j~��;?�"�` %Ch�#4��El�-ӭ�b�uT�K�ݭ��.Xc��k/�j�2���XĘ�R{�1�w��_&�??=t��XSƨ��6+z��먱�q�2�
_�$�1�(�M��qP�$B�u_��F�M�����XTi����Ow]�f��n���@ h0������rSؿ?"�� �[d�S.Ƨ<�;4{6P,.�~�h��a(#��P �L����L�¶���|��.=j[�3�P���.�Y�ڭQߑ�t�ʬ���T<��5sY�:�"oQk���Q`�g���+�?;�g�ۢ?���s�D[D<��9fѿ�̴^��i�<�r95)�ؘr��3òl������������a
$/�[G��g���
7�.��	�	^4L�h�G�2}�\��wậ��f�<m·�ёl��A�� Mp?#�MZ�SRl��Hj��ު���Ac��E��'?�R�֬Z

��Tr���1��-�O�x��E���5���v�4�p\��i��+U�@0���b����mA�ދ��D�r6~���ǿ��oX��b�+����ϥ���Pt<sjv�Gp���иƝU������<��4�1�oHN�#�;��J��	��-���z��Ȣ�	�kD�v���������W�i�na수�#OZ��)��g�H���e�dڡ1�P�i�J��8��<�G����!���3���;:=j���v�e�R��ݡ����Js&�Ýv:�����%=��t�(e\����&0�Y�������/c�:���SA}QvB��>@�ڳh��CF��\R{r��~=����:d����sn� ��ܬpb�;T1����OɗW��(�h�8�!ލ�DaU��+���tv��I�|�&�Ϗ�?]BshM��7��:���<hg����_�?"`n`�a^_�C;�ضx�� �3a�l$4zPzů��NO̬�-!�D���S[�o�k� ;c�;>/�"T��݈��K���ɟ������5ncm��@|�<U���6O��I���419_�-.n�����i�DUN��@m2�%|�Bj-�� ��9���ej����������:�R�#8��a��w^�V΋0i��DkQd4�B>�4�v2��*��27�n�*�?����p�ܲY?J�����h��`�歁����JZ;v�����V�}6�Õ�z�����M@�nj�[��n�/2zd�T_,�����x���3M�x�ȕR}_����KO��fY/�?ˎ��4�ߴ0�Aý����*�A.�| �/�'Y�M<YRq�7t���*�������
�|�p����K,%�8Q��ў}�Ѣ:�y���%	��&����+N-��F����l�P�]Z��
��(��7b����-r���T�2q���0{X��y�>����؊>���r0���ojWlO�'���1�9�����QED�c��$�IO�Bu��oV�?|��;������PT;����Ny�B��׋�$��)�7��i�1ֳ}�)B�����L:��7޽�2��1��@�0휯�?����<$��X���\rw|�+D������҆xN};(����!�"UX�������]�����=(Y��`�����G�E� ���Xuv��-�\�(�K~�����q�(d��y�\�q�M
��^K��0�%5�ȬW���(U�G��=��&����^�� M��m�D���a�߇a��*4�Q�x=�N�Zr4.�2?����7�ޞ���\���M��Ȇ�[�aD�٫�?`3�5�zB��D���k�om�ǋEt^P��~�9�PP~������Wm�X�>3�0���@�ղw��&��R'H|A�H�V���kS�Wo����zs'�*�^��Lg'��R �D;U��R���w�8??Y��8���
>�u6�RRsc�x����m�T�ѧI�f6b±�t�B� �z�W��i�")���ɜc�]�f-�6�s@I��Ǽ�e�mIc����[J

�|�F�y��I�l�.ХxP����EZ���;�sv^tro���)8G}f��E���2�O|8��ˤ��v��:\����}�����&y�͈��Y�	~k��>=��F/p��i�%�D f�X���s_}��:˔�,�d�wr���=��b���O� / ;rȴ�0X�֌��֦ŏ$��&��X慸�_?�'t�^&�Zs�f�����<b����8�\�-�f5�Wl2q��2(H��O
�o$ X�Ӽ\��q־�\�_U�pI0���x��6j�5$e>�����^���5���?Ԙ�3�a��{⛡��]SC��]�·�5����x�=�)l�P����ie�����zHOx�gAo��) ��������
u�IQ�L1U�9:
�
�^$Y�4�9�Y�h���6}�&��z��?�*��˴�8�F  �[��bX�hx ә�[���A5]`�ޚO�lc>��/ӱQ�^',�u��-���q�����,g��WTd����s�щvjҬ�7��}��O�|4So���a~�B��H�.�C\�q��~��d�+W]�tb�T�����@�Yn@�Oڟ���s|rK�a���;��37��<<��%s�������ҝ�[h�*�������j]��b�ІA�Zt����͛�m�2Cc�(Ȣ�=�Թ��KFY��3`�Hy�a8������'�xV��K���(Wڄ�jϐ�P�����1.~T��>VR,č(�kw"�,#��Q(�syqq�}qbo��4�l����V��Q5�TB6n��U�GΡ�P��
�ٓ��9$(�:s����Z��:*|#U�@.�uZ	��H�[��rz�{G�7��
u��\�jQ7k
?>fu� ��������TX���7�n7�@n�U�V�I�LN����?͛������BV�ȡ��HCй4��I�	�J��j[%��M�0���4l��c>��F4	wڢ�[/�(�J�jX�����q_]�j7�d[r��U=�I�Vl0�v�ݱ�?����`�d�"���ps	�N]U�j\/Z)�D �̹��>�"�DD�fP��A���$�-]��no�e�Hlüx |mr�a4�[ů1%wA���v�g�e�Ph�[S,��6r%�������R5��ͫUS_&ú�.K]�J8D�,ϕ=�U�g�)%A#���"L���QK�%ݸ_�V�i���0B`D������(�K+�w�9�����R�n�뇄�^n�-@�	�)�:��Vo���������Q�#u��cr��\����>�F��=����Y#&;����Z�	��pZ߁�	 HԹ+B�����C7#g:�h���}���=��k4�=�CdrX��K���3 پ�*�˞E7��#7��2[�/��&�|��O��O)=�\ˆ�O]�nn�*��u�����ΝLY9*�8�hޥB�7��fn"�V�h����y���	o��-4���s�H�t��[�څ��7w9�A�W=}�%_��E��w���g�z��Д~�Bb���#7��j-�_��q����n�Ǳ[?1ϊRP7
NM`z��٭)h�_�Ǔ2�"��}�n��a�n��;wa��-�3/���+%�w����b��u�}sC�����5xd3�V�\�Q��-��m��n�J������}%Ole&���lr�7��7��樔!� ʤ���.E�`�WԦ��^aθsUMl�=?(�װ,6�	J�%���<�B���?�WE>��<��lhl&�?���X�
o�[UUR
r�_�jnb�:���ݳO�<�����kN]��)��4��Cp_ݐ������:F�z��?tG�jh���s�>=�d
��T_�w^�}�>�FnċS��'�y:h��ӛm��z:���|0@$��&�M�ǛVUΜ5i���>y*��=��Vn�03�?OJ袭U�G����4s�!|� *b���l[o��W�H���7���: {Ұx RTA������6槽�iO��}u�/�d<o�rU�<̊my+�_�bn5��"㑷o`Tbl�81�mDP�L�8Ě��l��Ⲕ�4�[Y��>�{#�rj�'��0-A92�#;8S��<H�9�]��.�'_�H]���!XG3L��	S���L?/:�[(h[l��70�=����z��|�U�)��.*��%E���]}���e�h_(��3P)<���tQ/�_&$�����JR O��Cn�Ֆ�lyԙ�C�/S�hQ ���Æ��T{��f2ʑ<��!�t���vh>1$����v���ڦ2�v/sh��P������+��p[4/�=I�u�*_k]��V�o5��P�6eӤ�O�)<�oe	=��T��g�HY6���~?k��ӂ�Py��vy�uSV��[�q��&��Tef�֞����%5�	���P>���ITL�#T'?*E�~��m�B�w����}P��gơ�����C���N# ��m �"�?�8�F�}s1���s[�7ɿ��@i��ζ�N}�z��3�
�X_�7Nn���R9��W>l�u	s�bw�yQY��0��.��Y���'��t��q��Sw�!���-��m�����9ɔ1����B���><�TI`4�_���Cj� �P�Ej���`�v.��#<�u�VX�b�N�C<���K��O�}ұ��TL~�ͺ��÷&�gTB�ҥ�ߩq���u`D����6sIhQ/0��ʢJ�+��i.@r4��T�"���>�f�8���<���f�~���CM��߶�����vX˖�p���|ro�{x��O��ӏ�J��/,����S�@+�-`�R�޶��%+�՟�&� \zLYϫȻ�� ���z:�Y�l��� 
�����[En~ԋXH�Ħj�u'�6��e E𜠍~���&���O�β�Q�֚S�簢�(D�����y���Gx�VFNR�e/$�]����7Ν�>��?ˡ�b>~�6��b��D��(VY����rbj�WY��k3<�Jx�&���A��V^]����\�Z�i=.+W����'��"<QV[�^�	��+?$������ 㷀���b��'T(���'�Ķ�_��?��<���S�����I�8�p:�vR�Vɀ��fYF6��v��E�^B6����Vc�:J�BKS@;����c.�g��1H�4N�մ��.��ծa�P�E�%0��>9f'����x���l��;��hl�?�~G����7Ff�!({��1��}}Uȏ�P��� I~6���C�b�hR�Y���|���0$�$]��Դ�ٳF��ɖv���Ru�,�|}i��[./�SΤXe����c�6�U�a����<Z8�B�ƍV����;���c�_l;���06����[�>+C�]�I��=��iQye/�ĳA�A������o:`d�D�P}n��m_�vA�T�]��S&ͣl���"}�S��
ܰ�&e_���f�bO�t~�:V=���R;[]�8���U<�T(fԛ����*2GS�}�(/��ƎY`���}�;>\c�N�տ�yL7�<��p.�?��ʞ�������m^�+�!Ku����j�r!~�wVou���xL+�![𧫁Ƨ'�~�K3��A�O2H��C�u�r�k��ݥ��F�术���|�.sI���й9���7�G���qo)W��%�`��9���>�8��Z��Į�$�|}c�۾��`��ܿ���<��~X�������7�0w���g,�A�˙s�iİ6_Ο�{*�Y'���:�Ms^��_���+�^t���{i¼�9#����L�xj����b�k��*� &���Y����6��CCCF�{T�~r]���2��&���W�⫠φP�Q����J��E>��ݢ3�<7��L޽E���~iD�J&���s�/�������a������=��
S�M�G<bل��2��ئI�R�l�>s�#M*�N=�!����4oLI�Rh$(Ԥ��֨�߶O��4�������[������k"J���L*�IH�������E<��(��锇��z�Gf{��o�B'���eԧ%������lX+e�ח� ����/3 �1e%��p}����}�t��Y��y�Zl�}���%/G�2�m�ww}2�ii��"@�c�l�b&��8"��խ�^�/��Ʌ��`!�V��@��R�}�剆�ୱ�����5~@ՃG���X��zB/�2���K���)ء�2�d5'��x4�c`t�ڳ��B�����ů���]jN����l�\�
���.�?x	�5p��Tݥ 2������&SEf�ϛ�����������v�&�/���<]��\Z��ީ{���ֵ7tP3�&���� s���A�8��r��y_(~^{jk$�[��*sM��=J (���av/fy ����kO")ISj`��B��8��z��o�x�^�dVQ�­�z��h�� �ꗂh�]��{�h�%��t��9q}���?d�7(#ԇY6���|���}@��.�`��Ҝ�+Dt��Ռ`�1?"<�mj���r�8^~k�jb�"�*��}NW�߳�Ak��i��c1u6����s?1�^�-;�ia�畋�nݷ>��k��*�Ŕ����	&�&�)��m8���0�="�4���αd�C���C�E�
�RRQ��	=���<.-��"��f�9�����(��#����a;hj`�o+�<�ѵl܉$��Exs7T��j��ק#[�C�����B��Ȉ�3 �b����hLl˖�7�ͭ3����[�z�A�>��P��A��М��m��],�z�������������u��4��8���D�JQ��x}?4�>���k�H�T�H�_ǫ�V�^���؃��<v�t���͚>��!:`^s۴�k\F!��o�y��t&$��Vt�����^=�@uD���F�&�1��1�Ԓu�D@��ohq�{�q��P�W�8�I�=B,��"��{IӘ�b�
̀��sth(*%���Z;��S�1�oY+�OK�<-A'���O����j�x�����]/<����� �fh���Ee�ʏ"�����1k�w���p�D��@�b?�_ b�l_]����	�>��;U�29S:y�.s��:��zX���6�Y�eU���
�*'e������ň�����:�^u�:m*I1Sz�5cwԛ+Y?6'�9�(�EՍ�
�'�o�Xڝ[} ���`��p�2I.\lK�5�A�0�n���My7;�x�3���8���MI�h�$*�Xx'���0�U�E���4����ז��:�<}~e�}0xէ���%�=y˸b���^�d�7)��9�N8��������=C��=a�7@�v��2	�-���s@u3�70��GgS�v����z���@W�ҿ���
�2�YJu-Ayj�LT�����gִ�k-��@�%��g�>Z�qf� dt������k���t��J[^�"�&�:@8�c����7zjx�������+V'�[hLY17}%��nV����\`c�=[��7�)��x(H�8
�>GAų���F���j��AG]������N�9��9��Y��c�j����xJ��^P�n�MC��'KK	E[�8O�9it_iP��\?4�^�A5G��#�_����{*;��x(�57��3?[~��p<�f�2��|u��D_�颭TS�K/��]��S
��̑��;�)���lQ2a��~;h2n�Y\�T�_����7u�|cQ�	2���\�7b.x����/[�Ҁ��*8�_�y�9�P���{�V����c�ޯ?簀�#?��`�R���D�Ìޅt}�1���3�ߔ:�B���,o_?f�t�ڋ���.�F �V��ݣ�)�S?"��U>�+�oJ�#�O��0��.��,�wڊ��u���`���5�߹*�0yX�,�.-N��%�Ƽ������J�A�_�[�w�.���>��BAQӰ�t�������J��@6нZ�pr]�*�nX���yZ~m����G��F����س[�\J$��a�9>�#�`�)M�s~�����#,������o�=�ⶊ��ۘ�X2��op�sG"	EF�;�qz��rK%�⸗��a��"�d�\bky~GȒ��ÅSvw�U6��8��Q �E]��eAy�.�f��ք{��f����xi�/,���!��V�,!�.�t���:��6�*V�Hb�rߜ�S��+:_լƚ:�2��v9�imJG,�$����*� �Q�u'Y�����{M�W��ߡ������M��F�=ж�P���3n�ۤ��v�'�ӭ����>1 
�V��kx?ğ�����+�[�`$��e-�� ��M��
���HִޓD����W�d�]��n|���(���}u�x37�H��ZZZ��Ү�'�}![��q<P����~�q����e)>����Ħ��~���#L']���U��Ç���U������t:�aw�A�~8�U,�K������������PD�J�P�����N��I)	���B�%����`��=s����/_��f��{�u]�^kOQ׸��O�҂�,��I'�>�pR#ϕ������]�I��k"R�(���*ϑ���W�i����&��]��5U2e0�t����co�����;o�cպW|���#��Z!�_/Wa|>�[�X9�}��pYX����z|'t�ӄ��;�6�ٯ2������C�C�\F-���U�z���t�������	�2��{�m�^P��K�m��L����m����N&ǅ9 �梮����Z�I�)�#tx�̸� 8��;Jn�]��-�FX��6�q��2�iۥ�gf�a-%Y��^5z���*6|(�y��@���
,�������l��o�N�������n"�޵w�;�4v�߅��ku�9B�����m����޿a7����K��۵�gR�M��$�����
�m�Z-��]I��&�̏�ҡw��v�0=��4�I޷Õ�P�"覃�*�������l̤^��C��~��<N���b�;g�
E:��.\�y	��;\S����'~�d&%�dg$$G}�|:	K}��U'b<�k��I��mZ��W��
��m/Ե�*�|�[-�.���X?<�Zr�ԉy�g���������'�0"buI�͟K��b}�j,��0��Ph�,֖?"�^���������٨qoh����e�����z&�B�ߊ�#]�<-h����A*/��������Ii�����Ir�2m8ΐ�^�g����"����M~I��6��H�j����"�����V:�!�NF(���.��4�g����r�������+b	�:����`*ڸu}w-�u���? ��rK�U)Z�އW��U2��U3w��"+/�f�	\d����Jp���9�+�����L���R�StÈ��~��@Eb�l8�.Ht��߫��7�K�#�5�ɛ^�R�N1�B�����*<2'���3r
���H��5f�zL�	��t�;�k,(�w��<��S�ݛYx��+3蝞�|,8���vǆMLLLU�R�3���:X4@� zCy�Q|��x$�&#�(�:,�C�XCDI�wH�$�ff4g;^:��Q�S�B]�;WU�Fȹ�~8۪JJK���:D��)��׍��� Ϋ��K7 �|�ւ�lL������
1CH3�nm�g�� Z�'{���ힹ
⓾��^��8��Ǆ���k��4�� V�l2�@f�@�y	I	qx
����+�m��S��=��fb�n�/���x/��v�	������o/S%|��^#��7r`�X5��k}oZ���ەl�}밭i.dX��xR�E�g|����fY[u�}��!\u�qq��(�F�e���`u��qR3�]mp��(�/����M��Q��Zj��%_���i�Ηo�[�?zR�#�������%S�2�m[��_] .6�]�C���������*������[	��k�)���I��D@@Ւ���C��t�p��.�/�/).����T�� t�5D�vf����O�{���e3�fS��J�;��R+[y��%��:�dR72�{C�OWre��"^~�y-�2i�"^����k����$�AvG������&�
o���Ӈ�ZLn��^t�}�/��|��f�aW�F���?�oU	�.]X1�\ˣz�lɫ�v�2����)ߣA��h�3 L�i.f�kK`��j l������`[��!�d�u����3[lH���EW:��}=��%ȯq�(�?�g�U��`gozL��\�EZ� ��%#3��qq<�Weg�LL�ω�E��8����1E�r���.Z�]�	>�� �ؑ^��Ď{b�l���-&��7M�X��a�}l�f�R##�Pr�S��TM��]s.C��%LJfB��1gs,�E����LE�~M�3��.U��(�>54��n��з4����R���u�}����Yl��T�#��������g%���#�1�����d�I|n�܁�?�h�p�5�j;���.�h�7q�&�JzVgFFbg˾9����Y6�)5J�b����^����0QR[oc'KODi������OT�{����VR�<E0�����g�~�%J�x1�!�����rZa���~	"{�VF�45d4Ab�g��'	=u��ݽ�c�l�~>�Z�Wκ'����)�:;�7�L=J�|���R���Xg�e��]]���{�N��v^�%�zUJ�H� ���Q�w�"�y�7{w���;H�.�W�'��=D�������v��鐋���`���PP۽��?��c��O	�hE�j[�|e�Սg.c�<����*@��x�S��:!<W/� 9"��<�ιD���H�`��}k�zh �{�|A����͏�ﶡZ���J�����`±���3�8TV*�L9%#C
o΋}p�'��oN�`�(�u�����m��z�G�wF��6�+��y����J�����}�6�d�	�6���l���F�� A�i�쑚��ao;�B�s
�n��""�̼ U��xlMԴI�@+��8@���y"n�����z<9�4".�񝨈�p�3��~��YG��ָSz��d�>"LJ�$X�|!��$�P0k� ��g��C}ڏ�@�U6���y*#�o� �3Ԯ�MZ<��<wR9��e��%��&(���j�I������>}Ї!B��T@���;r�HQ� 2�K�4��C�\�_��Zd��Ej��^�mƦ����7��-��|�c��`��V�i�M����B?�r7R^��0�މP��M��K2;n>ے,:e�~�:LZs?��_�M�$���{"疏
t
�j�f�������	��qu��GF��)����?��>����F��2Ui� � 5_����yE͗z����� Ȝڸ�+����'��Y��mX8�	ȏ��3�!�c���G��j�2��'<OʡXlЌĜK����̴\�r:ǑS岯P�7S���KK�u���^`�m۝>����� �9�a�Y�uYr�������AOh�Go`\m^1�y�1�[��j��H�l6�Ug���Bl=Ja�4&�����f^���r0���1�%%�40x+���Y0�W�_��П���c)�}���'��,��ƚy~����7K-���4�|�{!�u�	M.b!�%!��F~b�H?U�{\�"������m"$edB�E��4���G���<�)<j[��x��i@[@�6}x��8X�(E�6ӲL��낐��͇�4�:@��-RS��A�2����]}oNY�x��$߯��n#�]*ܕ-A�B	���6�ˮ���>#���S���/�N����8���U<c��?(�Z�oM�7F�GƹSf��g��f6�R �Ȱ&0�� |��\�ǝ�y��ͅw`�3�DƂ��;�)�3T���?Z�ѫε:�p6����3�p��hAQ�����>�_��21��w)�?�X���N���{�;~��3��P�f
�B�1XO��Id��n�i��)�i�����58͵��, �j�*t{���m1{A����9��|i�/��rzY�أ��=��k�6�2/*��˕��^!-�w_a���6�#wW���]��� �����
ᜯ������.wx/��<Ż�u��i��ϋ�pM�`�U�#�z4>�^��490tV �H&LHL���y��o�eT���B0�iVT�[CQ��'V�u���-O#yDȋW��Wх��B�x�2z (�Oo�V�6�?���|�0Zd{�]~7�is�  �s"(�/��z��Z�h��7A��o��� �rB�Z+m�&�����ߎ�^Żˤ��u>�X�v1�D�oؠ����,���E~62e;��ì3;��.�,�k;��`ZɁН!	�y ���]qv ���.g����5�c��+W�R�O��0t���Ӱƃ*������Oe{hr>ʊ���-^Y�5�����J��Z��}�u��P޺�ZJ���N����A����7ؒ]��%M}b���Tu[M`���D���V�e�X�Ӹ�x/�)���s�f�u�V���˔�w_�s4�'`z	���ckc�v`�.暿��j��[�{ە�<&$�
���AdwL;�tGw��`'�^ʊ��<��/���u�B�(w�L����M�&j��dj���v>�7-c*i'��pO��egZq	B�����62���ŇY�ΰL�(�e��K����[�&Iqx]
c�F0%�ț ��X~�b�"׋�U�a~���X���x�'��^"����{>%���4 nAKy�) |0���5�n�c]�М��Y����ֺ!b��{�m�Q�/}J��#��m!�|ݟp��y�=c�#1m�I)�?��n�����r)�2>��-���w�k�/���=w2�d˨�����uS�����@�Q�U����b�Vp:�zp����^VX,�h�r�xTㅐ��~��P��WNug~N �đ�<'E�C{���o�%�w�K���:��7�rH-�4XV��F�����49�^+f�Ln��Tx�������ab�Ψ��ه���SV ����>W�;��8e�g�0��e�E�Q���WRH>8ht��	�b3���}���g��O�o%�l�Gا��L�O�Y1�W��V�#R�/��U�˱�+E�CJNuz>ƎKį<�^��te4��}TKk	��� [��˘z��dGү���s_`N}ًD�;-�3J��-UU_�k��o����R4���-';����,�W�jc窄wb
}VK�I�J� M�/z�*�H�䂖
-���A)j5�H,~����O��h?��[�[ ����$Z�V��Nf����4��Sfv�e��8�-�S�1{���Ib���=[x;?$�fZ"���̙Jơc=���ɨ��i�Ѱ����r���U�����î������´��^�������ߥ�*��~TP��6�|�H/�zF�LTk�����=ȷ�-�ZYn+�cqb���J��q�䏻�����;u� IBMVG�l���*M�J��Ċ�"hsC�2b���.�T�(��|$LJRfA�J]�ׄ�_V��� �[�Sj@oU�b�9����ӧʂ�*̳u�I�D�5����("3�{�����=�1���Pi��|�i����dɉ�
l����%�	�R�A�*=3s�i�L4R�Wi�^�IQE�F�V^M������Z��5#�e���q��g<Bs{��܋ˮ�o�eޏ+��VW�W�>�ݥ?�k��߷���"��l��8�o�u|9f�3�M6$Y�*��QA7ݶCw��0uE��ֳ Q�3�6����C�&{w�E"����؃����y�L����UY�>.�����v�
�"T����`�m,C�%�4��AX�`@"��{R+�)���i�W�1g4�j1�_3�1@���J?�����'���G��l����M�w9����um.gݔc�D��w�h�5e��4D��5�x����H�+��7�Wb� �Q�f?�z�֚0�5�}jں�������9t�m�c�ζs���L~�[�$^E4����	�lL�K�d����{�V7XФt�4�����"�bΤ�����Z�ʥ����^�g�fl��=s��*_�l�߯����D���!%A1ؕ_�Ɍ�n��`�_�ǯ{B�_�Ní�{�C_N��q ��^�{����v-� ����l��꠼�uG<��	%7�� N`'	7p��&�C/��J"�;@%�W#oZ�_��O���юU�͚I}8FS��{�[Mk�P>��{~��uzPr��m[o�n�H�wH��!c:����~K;��AZ���TѴ"ޏQA�E5S������a�էu���i�5��]D�dS�El�b6�%\º,����)Vu��@,s붖_� ��J���O�$#���W!�H�:�Q�f�{�l61��:#e���i�L���x�¨*�w%�}Z��xl<�ɾj	��1�R�
#�ں��;<�"� <F�V���d�O��V6���U4��C$IeG.(�D��I�]�Q��?u�L�D���2J��w�tyKV
YflؗE?�M|�#s�ސÛ0�y+ѯ@Qx��ҋ��3�kO��>d�@ъ���?��~�U�i�O�{9��f�X��Ղ.��<��h�cĘ�:�| �"��xFR��N����� f���(����pbT�����Ҩ�+��9�Cu�R�[�gbj�˦�G`Glw2��ot�'��&s�֞��Ҙ����1Yi@Td*����$J	՜�)�MD�p���HI��պ�df� ��E%>�S<�ϗͼ[�˰� �eRl���;<�� ^~X*9;eNE=������7n8��o����H�Fϗ�	������A����z׆���lHN�1�������R��r�8}?/�N3����u�ݰ����r�Ʋ�g���+����;�J������׉�Mx���ð��+0��!�l��qsp�oX��+"�|�/rC>�Edn'�F�������6t���?fk1��}����9[�H�e[ۅ9`qThx8��;Y�}W� �&���w�Ղ�	�?�V쪴h��Gx��匊*����QXT2ELy5W��69�R�])�_�9�H�z<��551s�0T�X��������s�	d�����)%to���+b:Z��&[������\a|��gEx֨�����|R���s�%�_տ�`��<������+q�4u���Bf�[i:��NX�efW�vm-�=w�xC+��H|8B�5�iL ۆ��[5��>P\�#0(�$�|���Y���8)�vWfX�Z{9u%����ږ�����UF��w��l�����~v;�}E��]a?�Z����cP��#V#}��]�h�i�\��5�kcN���A�0�Jv���h�`��2���@�PL�}�����RsocM`H ��שː���O�g���X.y���
b�B�=�Z//�Q��'�٫�UP�)T������gQ"�}Et�=��!a}SJ��x�%�a�)F��L��J[G�����h�T2?��
�#^s'{��6�$�S�[���Pz���&�y�K���I��-��[`L��틁�~�	9Lg>����21-�.8��cj������������lB7kKP���\aJ���Y�	־m���_{��o��R���yq�a[JwC�`��b�����Q�GL Ď�gY	�$(B���s
��8̆�(�?��NH�):{y�
�x������d��-E�&�S���G�̩d���v��oa����"���dv�w
�l8��\��\�� ]�;:�A���y��Ұ������g��n���$�v���xk�W0} ��/�uE���
+4Eoy��KT��b�zO��s�ލ3�ڳ���CŢ�>m6FC�6���d�ؾ��	�Վ�FmEm��Sc����
B*�A��Uw��W�wET�9����۶R�! {�7�vG̦0c��%?���^����ɟ���^x�%�߿THo��f<`���ᵺ�8�������ھ��V����/vph���f�(sJ�h������r�r�1I�[&����R2��Q���֑6B��ȟ'[Y��sK�^>��>?��D��WF�yh��WU&M..�� \fd�:�	�p�����s������I:N�0�~��%�28#�z�O�/٣�)X�47�Ccw���v� ��cސ3s<Sެ�����Db�%g�.e9@B��u�Wc% ��ս檆s	V_����gb,���%���F��*��2~˯��ooM��rNx�٩cJ�[E)�*]����g�~?��yʝ`�\w�+G��o�l�/8�e%��
Ӆ�"�x��ڐK;����j ����|�C�q7E������]L�%L`�ow�9��/_c˅�=f����Jq�hun����8]��OlM�L�뽹��$��$X��V�4N�╢��S��53,�x�g���)��X��~��v0&���9�2��t�pi}�'0�C1qVVF�b���_�Rb֏d��5�iY��z�喛��1�8��=o������җ��I͸��Ғ[uE0f?K7I���#��R6�����d��������`N~Q��;�7�¾�G�\f$�s��s���R���'��8�;�U�����/���9����ƭ�[����f1�}��W?ό:T��Wޑ�ɰ,-{/�9���7����J�ʼ&�'"�b��C~1h}�X�> �%0���ۊ��Q�y�(W[�AC�ݩEv�I���vث��o�7%����g���n�O����Y</�?�
�MG��7jQ�z��GM�~���A���	���������V��S���1��
���s�rVA����f�JZ,�z�x�������D�����&A��.���: ��-��BE�5y�̔�9�q=9��6�6�o��EE���5N�\U�jo�˱r��t����Fqx�l�$��OZ��3H�oU������jz%;M�;k�5���u��l֩�����tXQ��!�_5mx|�.av�Z���0�s2���&��;���=�ɭ��k߀�1b����b��}��~�D�²�Ϟ�<�se������Ax`Uq�p�x�b㹇�a��J9*p�������b�K߳�|c���+"F�'�� ���"Rxk�e#�D��(9Z�3�_>�v�3̢�>-�<~��LCyN�Bo�h���h6m<0BW&o7oX�%¨��m�@�'L�>=z�)5M���ߪ���=�Q��|;�U�(X�o���{S�^(�w�%�K$���]Z@�����1>�m�t���|%p����i�j��1�KS��o/*�ɯ���9,-�x����7�;�8�Z�e��	��i�K�9�n/�<�%ޮ7-�n���~����8�ᬪ�RyQ�?�����mT� W@XVRXA ^�@,п$�=[	�����o��+�N���>�'����O�w�����*�?
���b@BL���nO![X�_�����F��Ҟ��G��￀6�W��7]�fcSPZ!�>̭��[�
)���PK   �YzX؞�~O7  )8  /   images/ea12a0eb-7632-4157-afc7-05122dfed1cd.png={x\]�vl;il�n�4��8il�v����&��ƶ��i����:�33{�����	W��D�ÃA��&����Y��Ձۿ���QIR�r������W��X�CȏsX�o��  hN���k�Dn  \�Rb_U��N3��T������]�i������~p��A�Y��GD,�HGU�AF�Q��/����ȩ����#����;շ������
lL�oD�o��_K��[u4�8��O2&�677���R8��t�BX!�;��MKKk<��s�M4x9@Ĕ��7Q��΅�����=�g�F�Ʋ��ɊITZZ���?W�~��%�n����[J���*����6����%�pc;�����x�@SMM���}���&n�h�<h�laMR�C����:�@:u�~ݷ�7�Q���"��m���z�,U��qtt4)#�A�Б��u���aS[�Js2j���T���1�	��]!kw$uD^��7�$��Δ�_[��#~d���Ĕ�1�q�{���D��;xe��U5^SSd?R"^�p@�����z���Bh����JP^8�8K��S�l�EYYiA����7�rz���[,��1�n�K�?8�w	����
j|��l���^��9W��u��@����
�U��x8������V�W��']F�g��cTG"dӤdb���j�߶%�	��@�������'1	2�V��X�^�5k��3]+�5�ש4������s���&s���sK��¢���B�lKL�@rwBr:��qhs�	R���[>��LCD(�t�9���:j���xI�7�k�o�芘s��foe_��v���b�.�J��(+��QjX'V��^�7b&�q=󪈦r��J���)�.T���߷�<�KHN/�N�m�~sI�������:`��"O4�I�gW�q�Z��`�!##ӝ�}�P˴�3�	(�z��Q�$(0Q���L#4����ب����zq��"��*n�!*&KI�AV�χr�s���􏗡D;#LI���I�t�Hc�q4���2		�8�edĝlZ��)9�E�lj�o�*�*��QM	(ӱ�]�q�썦;���ny;F��Ő�54T�l�-X�x�A	VV��Г�!�G�H	�Lt��Bn�Y�3W�˶C	������c��C��-D!8��#��I�ô��W�����(9�H	�������$J,Ja5���[k6�k��h%F�&�,�?rk؆��~ЪI�6��0%t��d����k�t"MPԦ�TM���xi�ĥ��Ez�<i�L�TZ14�}c��r�;��6�Ua���nC��)����`j�Y���AYw�B	R����29<-�M�aY�1�M`K�#&�O��ŀߞ�c�2<�3�ŧ@d
�ӄ����o����S���a�-��}�*/����
ԃ�<)��)UTU�~�����ˇ �����G��Ư��Ґ�^@z}p��nS��y��H��W�|�W��K���j��I'%X8;mr��Y�t��:���c���[��݁k~�9�.�c�2��|��{�ܶiػ��M��њILߺ�3�P�g�i��D�
�	!h��V�oҔ6{=�+"�Ȉv(�	�eᲠ�Cn�~���2��JD�d��$���V�ȩT���P{?��[U��� hi��ڈJ�a-X�k'v�����^�B�5-�F4��L�.��~�+-+s�vJ#��#m�r/��s���*��r��8k���D� ,d�e-���6� V��t�*W	R�㑟�>E��������y!���\hAG���H�Ї�_�qI*9�����*��(��mm���U���d�����a���J{N)�!A.�j�����"��z<k=W���Bc@�x�*/�N�"\}���*�*@�l��#�E�x:��T�6GbJ�r��l"�8���y ���ܗ�9
�����l��>�������J�/�tTw�ѯl��g��A@� ��Iu�8hW������١�aK�q��2\!���>,�U��0	���3*Qp���T��#��n�m�M5U�(��r>��Up���H�8���5E���
�K�+5=����������2�xXNW�J���m�p pW��_�wO���O�낄aIKG�E/��i!��	M[*���fd��B�I�uX�<�ר��hv��[��0cE���k��R�CLbb�L9�d�˙��Zp&b��U��F��p����N^8����1q�A�P�Џ\�9m��a�ڨSJN�2)9��E��ѡƙ�R*�˰!�����%�v<�0��,k����>��p6^P�I���>�)��g|!��֟�vC��oQ��|\�N(�d�@57�?��Sc�9��j����6�G�DX����V�2@�����i~�I�k|���$*>0m��.������i4T�V��"� 9$�k���a���+��x5��Ǧ�_D�0Ȟt�X3����;�]E��n�	kT��	�h�i�������j�W!�5$�!��Q&��/��tH��f�}5U͓0��!+��F޾F�5p�R����K�q֧w���n�)U2qڹ��x�jX��kފ�3�#���ldTRcG	Q���Ӷm���:��a������b�_�2��25ߦhǶ�9�D������Hք^Y9#{�LI����&�,B�/hn:�O6o����ʶ��z���ߎdj��ނJ3�E01�1�[� �m>O}a�tn�I�R&�7gݒ^J�nZ%���b�����w�9���O�/��s�)	��/����� ����}d����x���\�y�-V�%�|��D���2��yڄn���������b�P�e'�����z�;�r]q/:i����@|1S1�EO�G� b��~��C� T�M(g�c-xEh���e;�\]�0��v�G��c V�y��{��B%E?���l\��o>�Z:t	<)���g$p�\a��}�-�]8��/��q�X"���U�rέ/�.��e���3~Ӣ�'�Sŵ���Ȭ�j�0�r��a�	o����=x�2����F>�?�V�Y��	P#X�Ma�;%�Ek�u$��?F�c%���-�I�[�*ŋ��5窛�*3L/�������W���(J�|�=�.�7���jrDE�0*�7bۤ��"e�7-xk�]��uG�+�xh���e��L�mG����8��-W{��o4u�g���P�D���v ��5̩@�Y�vvvv����۠aK>|��;����i���1�E(�����542h�u���}k��A�3F8�8�<��ጙ�s���AH���gIP��L�}����?h��b�qq�Il&b����[�v�Z�FC�{K
-�K�S�,��xLp���|	�}B��*�x����c����w~"�MhKMC��fK���9�Z�Q��  �LSp>[���߇�v޾JC�\���I��1�Ԛh��(a1j�$[�zuh�������7�B]���Z։��>�M_ה篦��T��W� ��e.�))ٮ��Z[ka�;.y��@|��H�Y�Ul�64�7N�Y�R����ˡ�kgۜ�#�Ĉ&��N���	��ܯAUP�=�����Gs���Ys<�{_4k��1*irKJ"g�4ڤQ+K��J��h��Q���î�ʪv�m;�?�O��>x(
#6Ӓ�1�"!��3vّ���T�yq��I7ˊw�B)!�Q8i�hA�B���C2+5�y\�j,��J �Vٗ9�����048<��L�/><�+�N�
t�j������4ו�,{.;@���'��#P�I��R�[���%~>�54�=����i3��ꎖf�&a�����Ŷˠq4�H��ۖ�L"&N��} ��e��N",~5D�=XV�N;!�^���t���H�N�� �n��y���@��&ZB�i���@y������F*�����9T����&�!��_�WU(�����nԏ�~�4�w$��}k���U��i�-Y�)�u!U�|��ˇ4�{ 3	�'���}�s���w�c������	׼��5@��{��D��&��H��H^k�������ԡ��W���E-LA�Fm-���ǧ2qV������TW���At���<�A�&]��uD��"��v�C�bd�U1;_�+� ��S=2�4c���m�W"���߿�p#(�}kV]��b�V�)FL�TǓێ��m�i��E�7�`�=P�6婓;^Fy@ɿY�O��o[�G�+�GX"�����vY~�{]t�h������ n���<���c��%��z]�d�h/�nWc��z;\sGఅ���J�i0vM
՘�"]b��W�bx��W�N��5œiNy'��egA!��GyD� ^g��^�57Q9�G���� �p���0�emgWآq���%���`z����
OD��<�*�����<������`8
K:���8��S���N���ޱk���9�z�\$7�7�~�Wr�uuB_,YE�-/|8��� �Į��E^�Am����a0��$��=�;K��w˶��ɗ�?9��y��7���2�b�p�5����\׽+W��D*�x�ۅ弾A�K���c``|�����>ʹ/ԏ�r	d��J����gOǻy�L)����cT�+zN߿���U��}��ǅ4&᳘�s���
d������R'�c1�"[���춤��|}�����N7U�3�e&V�z�����Jm�r��v=������8��:*)�nb����JUj.w���R'x�9��h��v�ߟRu�o�X}���!����dk*��� ����9�Yگ*��^? ���c�ݒ�]�C�2��}�r=�����դ(�I(~ V@m]��<~^����"���z1��c�Q�4q��2찠 ݙ~�Uk��ʇo�b�S�����3�,�L��&�/0�?�u��>�p]#A���p�?����z�xdm~�Nr%ߨ��cj�2j���m?:I7�4z�nw-M���5��0�Q=z� ��1��M���s�T<\��%l��6[���E��B��!It�g�(����wU��P"GL,f���v��긢a>�d�kɜLU���5�ݽ���m�GH_�}W��b��q︪v�kGŨ'�a�-{,�O}l;�:�sS��4����/Z���VE
J&�7Zj��~{'/�QɑX����V�ũd��#�q���3͌Вt�'%�G������zG�Pet��^�t���uS^��e�k�7�DY����+�	�z �k�{���Ⓙ�o�P��@�<X��iy2���p�_jF�x�e��m��Q3�w1^(b����M�h�£#�.��_��٠j�z߁|��^NČ"�f�ޔ��.�iq?<\[���#��(&.�&.�M����I��T�N ���j��o9�\l��qC!_{���K���y�۸��3<+3��iR��n��Gwz�XHVtC�b��>"�"Τ4X���B�L����e)�B�ew┭�P�(hʇٕ����d���oO�[�3A�RJ�fz%�|�r�UG�@W`c�Ue��݊�<-}R�Y�4�N��Kl�~և���B57���?�>$%�XP��r��jչQ�X/��-q�R7���NҞ�����gɦ��e�]���pw(���iQt&UGx�e0�^Ŕ@�l|�/�GT�n	'�A��Q2%�?r'r��2�3�1���U���OB;([1Bm�JbOk/�����Gq"G���	JZp_*j�����v������|����>��hp��T�����&֥��0 �Ͻ����2�����~e�/�t	�����1�R$��eJ��(�+զ��8-����'x�t̻�?����5�!�;EۆKP��ߛH%tS(��L�+���S�őm�<����T,`jF}�黎����Ѧ���׷�_;;ơ{�]��(w�
(`���G�ۼ2Z(Z(O>�#����d��IY3��L��+LV�ir�׺�k!g1~%_��!�L�s�7�/}����MNF�[���K"�. �Il�#�0iR�JSO:<�q��GN�iS��g^��9D�0!pPiْ��@)��I��!jE�"SO����uHD���r괒W�f��6˺W�xJF ��H~-����MҴ�H�N��I�J�:,&�.1o��UJ�Lfh=o�}�x�pX�����_(������R�a�vڶ_	��E1Ll�@~�Q��N�$
Խ>�/ԓ�N�B��p��Ԕ�\�IQ�^CR. ��	� nQv.�==��r��6c���*�m�m�m���fF~�Ȫr~�4حQj �&yi�Q�nD����@�a	2k4B�OЫ��r����x��/=�;o};�J}��/I'�F�嬰�������H��:�s@�#��?����������.3�\�s|���KF�5�|����_�Zm\�� ���b��q���|^?6}��<�i8��I��_�WQ�=����U&�B�f��HQ��'�%��FM�_U�F�o���1��Fap�MU�M�}��m};(��Έ�iw~@�W����LS-W�X���_=I�I�=�
���d�<�;4}Ϟ)���c,Q����r�X�:�ի�ڌ7:�y��H)��:.C^z��y�q�r�f?��4G )���?�&v��P�T���ߡ��Qb�1Dk ,����οh�B!N;�s�/��gK�Ӊ��Z���2ڔx��g�/t��.s��\4=�0���kʨa�����l�X�5w��2.�v!����t
۞ވ��,I�a(�A��>xF���D�2wR��^$�X��;JE����7 �{�M��[�v��nP;�_Ӳ�LVTjj����D\&9�D�(��]Z ��v���Ȇ�*����J�#6��H �A��`'^�K$m����9_��WcS�>�'A�a�?�������
܋f�ۧ���MY��P<:� j�
�[T��#8� �$���ob�9��_NGҏ�+~"���F`��_O8C����s�`Ĕ#PNBRݢ ����j��WV������+���_>��� m"<��	�3Փi5�nk2̕��-\c��ja�34
Lc�Qm��	A�, �^���d� `p�0���<5],Axɗ��~��P *���j�JS(e��� - l�Q+��r�XdS�%~�ӗ#��PlVGE�{�O��kW[�̽4�D�?14�
�t4+5���Tq�o?�@&�+�m���GQb�4����0�EE����	���VQm��� �
�<�2�c�*l#bNwOP#%c&��9Ȏ9G	ߜL�B����jRd�\#�.u�ݨ�a�,��y�,��~l���.#;�<i"�%8�7��-ɘ?e�YN�`2+eI�h������ЄLF�wa32)1�v_�O41Q����b^ ^0�dm�Jؚ��j��g<����BE��_���D�0��?f�6�X�y4
f���G�x�kX"\�*�Qf�����SPN@sD��;p1>uA��/,�����(ٰ�ښMcz� �O�ը��N�i�	�c&���p~S������Y���-�I�K7/�2��i]⸔�.���~�3���a�I��`<�j:�hiZ�W]#��J�ʅ�yP��\��
T7�=��r�jRY�aP8�Ӄ=�?81wou��2>f��I�(u��9��׈�x=gzf!�lt��_���%��L�a @��\���c!Kx�_�:��}�M�����b�7�v����o�Hz�*���b��y��bި�:t�ۺ� �}�<ng��%���@ōu]U������le51�� ���[�|!l���À	��Ă����E�r��Y4�M���cS�lq:-x�Ͱ{esEpm䦾x�w��S��#K����-��� (B�!+q�+���4��w�B�J���X���s�;sJ4o?��V5h��n>lv��31$�\`t]����$�u�GhzR@�$��* �����{H�~p����zh�O����B74 �_їE�a�E;�{8�����8Ę���K��Wl���թX��l7)&��g~�u���ߚ[5m�X����� W�̷ٔVk&��
mNVnw<� ,����3@�ϖ+b����j��p�%E5$���z��C ��ؼ�v���l6�F�E��L�U�X�.̭0{��zo�%�B�]��7�����n8�`?�1F�m3���d�ez7d8]M�yr�hm/m�Gbe��J�&u-[�i۶E�@ԣ{��Ӭym%5v7��Q�$X��N�&���N"
Z;���oPV��C��0�qH"Z��Y�5��5#6��9�
���2�+^��U�W�;9�>�:�/��\C�\��6m�j�v'��	�	��d��J_�v�	���{��Q�\ oG!�Lt�YE�5'��S��_�d��eO�j+�?�%���6c*]U�Ҹ�1��d�Ş85�<�e�/�j,�a�Cri��Ȑ�n:����K4^��7�L@b��6kX��뤙h����Ŋ�|�����"�ˈ��â���ks��D� �'#Ę����[\M��EL8���B�]L�@�@�������*f���:��7�Ś�ֆX+8[�`� �N���n�(R|�4�&���`��Q)]j�{f�:��e�*g��U��j61��И��r�V_�΀��r&?ݨ����&��^�A������͞��Fuwy�lU�A]�F&X��N��z1%Rɧܯ���@���x��1�	�a�%�l4�;	Hh��L��Vڔ���@��D[}ƃ����{�x쯷�ȫ�DyK>c��L�l���A4���\ _�[��'rv�9vүL]oE�����fw��5[���$Gz�QWA���e��:X�G�=h�h8Z6e��������s*�tܫlu�d)eʑ� �n˭rƘ
W5�ʝ���-/�*<��Y�Pi)Ŷy7�v�g��ǹ%�D��P�TaÁyv�:��-'
�MB��=�u=y��7-�6 �le\�Г�;ƣ�N�9�����b{�y �g|no�+P���gݔ���R�ݦ�f�Ӕ�hɁ1��-�t`�H�Կj��R�\�kkX�u]��l��+���3·�@VD{E��POSqw����X6_��B�筚q(Nw���[�o����6�����}�9�A�S�*��q$D� �{T^�h�Ⱥ��a��֟x�ʹ{�b�$8HQR�����P��o��o�'2���.�v���Ig�-�΀�W�l��l�_l[�_�;T��I�$`nLR�M�U�!!MzQ�i�����Ľ�&�61��/��Ĥu��
�L��ܶ����,~ܧs�Ti���ݠ���K���>��z{ܧb��I��JN&��	��R<�k��� OB?�nk�=�aZG��F1K��A,;r�g�]�ʤ�"�_��E�cSN��y��5���/K�`ŋ�5��N}�O1�qng��x	��v��K�Q	2@����=/��Wn�zWM��� n,�D&��|y\F�1���l��h/� ��^Eߤ�8��~�M��	�JD��JR�S�'c8B�CYqY6rM�� ?�
�GW�n�ch��d����K[�f�o�����z�@@x�����}ܫ�!�h�]R�MI&������	Gv'��l�&[�ޅ^�Iܦ�%����v�j3I��n��\�~�t[)�/S�t{L��9֒��VA�T0�z���k��W"�a�_�~�j�Q{��-�1WN|�wH}9a���(5��.談�ؑ��g�?4�|�\���(n>1�D�:,��UO�����9�-H'������>Ѩ}޹�������D�	�|Z�|���$غ�T}M�j<\�)�y ��˟B9�[�OS�o�V��Nb�yL�>�g��E8�:��!�c���Y�M�+SD���(��W���F�����@��!�Q�����d���O>���jz�Q�>Y5?$H/�6�R�wA%x��J�v�.�I<�с=�7����D<��FF�Yh���R��-$��V�"lN�����R�ǡ�n��YA�/��|����o\	�[��O��m'о ��1��L���-�#����t;&^�E���D���kD'���k�]!���]I��~�CsW�&e���8�5���V F�{e�%�Xv��&�4�ð�<qֽ��l��FE��fz��K4�$*��µ��� ��(��L_�)Z���"�{�!�2��)���ZE��Ta��-����j�m鳶�"K�y��(�W7�A++��(z���ւ`��i�jxU���uLG����G�K����r���a�u�yy:�sc�2=T9�ަ�dg��?���~�����	�x2���s���e�)�����i*R�S�t�4�(��P��
���˘FKR�Ѵ��q@��<���;�}��8[��dU��v���9y��Wb��cɡ�'|N����Y����T`��k��t�q+�)���5xM�0�C��u��~b.ٕ3���e`P��ņ�ˆ_�q��w�U�F	��
�B� ϩ#3ddiizm��ƣII��VH%u�� p]舞��1l3-s^�pn�@e���_rG��	���P��T7���Z���u�ȗ�3gvC�|/=�h ?�N���PQQ+>T!F�DC����C^�τ�<0��`�dG��@r�+�+��!��R �͇�n�Z��tD�*��C�|��ݬ��=�=�Kͮ�-"�q?�����&|p[�>jr���("\<��d!�XN���J��RAᏒ$âYi�[�h?t%8DD�yg�w�[�Z�}3����|�(�I�z�����J�0ao���Srq���<��FA�ä4��i�ɩ�U��d���iz�@^{]9,�J���w�K����I���Ӛ4ͷEȪ��N�M��(?Z�3|����%;+�woz�c�3��y^=�oA���z�k#+��g=/UtM�F����"F�z9D�T]�h�>��߼��0V|�>k�"���k��N��ʥY�I����Ri\�N���7�A�'�?iI�ճ�v�j��<+3���s=�������bN+����\��Q�K��VC��YyO3�Iq]w�j��t1B��KظbI��J��'���w��X�܁�OdME�QߡE���"Thp�D�9�j�
�jO�����_�	f����>�s]p��6哷9�7K!W�^��ϤE�+�����������m��?%����������9����Ϗ^�MN^y�t|�eX�2%�'DJ��?D�X�#ǿ	����P����_vO�7 {�I*��4�r����ۍw;8�����yt�z�R����4�=m!+�K-ε�"��f�lݨ��/�qc4/��B"12��<�5$;K1�%���*P=?�q����$�]��m���j�T7��^�I<Z��v/��|ޡ�j��!2�y��c�ua2�x�	n|�� �?��uJ1���1����SՒ3����܂��7��V�;X
}��-^�<��ir*�C�Xْ���1�N���~���d��9��`CXU�r��W��x4��+�9�y�e)W�u���Bs�I\H�A.22]>��Q����JSn<��O�O�}�d�~v�a�[u\ա���O���E �W�'���-U�P��`tM�+�?����uZ���k4����,�鿅��zN�Yb"�@x0���g��=�|_�}��5�	��T��#�1.�a�{�H�������:*4ot�;��[�T�I���흓�7V]e3'9,IO��A��Z�&�'��J�D������Ն��(w�~�_0��wx_��~Q��8�ߜ��W����!���;U\Z���ZR�FҸ���rу\���Us�d�:P�I�zZ�_`�p���j#"�+U�|��?�3�����q�}��(f�V�mVKt
��'�s���q�41������_�>N�zN˝]�sf�;Wο������#WT{�5o���7�N(btl+-��uq�s<,�U�=F������\�C�5�E�c��a�W��aS�K=-5�"� 	ohN3�*�ˠ_G(���}��Mm�ŹBv>���J���V0����r�?l�۝�HI㏏V�SN.:�{A�S��>�P�����s`z~��$���J���C��W�O�ZnhV� N�|�G��y��$;�P%2�<	�̽�U�=�[�>��*��Oy>9�K��C<"LE�|�9;V�w~AQ	,���W��I��NL,Se�X��o�yanJ�	�d�byNn��C7%;4a�swZ���*J�~�]�a��dep�%h��G??��|��Z�/��bB�����x�m+)�����؜���tBۖ��O�G�?K��7�+
��|��#���B�|Oe7cV�]��P���e��C�з\� 7�"�o�4(���DiR���`Fhmi-����Y�\�(M�Z�%X�ʛ��0��˻���v�pɧ�*_�����2���΁Rr�����k�w7�k\��q'����L�J3Z'�H�� �+�YL�^�\���Ǻ�����+uh<�fM0��N�����Zq��������XK���k�Ȝ=\g��e�ω��*������I�D��4#�7t�0����ܣjZ��c�߆g�#�p����31bī�	(�J��J/d7e�9_�7~�2������j�	��V����ۙ�K��4�F��ƨ�%�r�fӾ��.ԝ�Z����]|h4�鉨�@ ��t�����V��{��!s������IѡD߲��`5����'�+��<�"�,H
��B��$���"�*�?����)�x0y��n�W�Dǯ�/��ǘ�cP>�@Bo��Z��y۷��0Icg|[jd[��z����;�TTÐ�n�'���ݥڶ�"���a�)��m�dC�=1�s� �ջ�>���#J&�
w5���J�Sa���n���k�x��.c}JW�򾏌N6����%�A�OH���Y�����o�w��Q"�C���x���C�� 	����c��6D �p������J�/,%��i!�Y�S��|��[�ccsF�&=��tB�-�Dk�����ߧ���B4����N��+1GR�/-U�PΜ�#L������(�\3�2ib�	!Ői._'�
&��5pm�J�e��E]Zr��Z�y���8*)4��*U-����I�g��ԩ5��/��ٟ.�h%��X��i���}���9�
`��@B�T@��{P�鯾��T�^��qRd,�}7=���f
��c�:�w�Ȣ��QNYH�CLFRJ������='��P�ic��5�ǆ1y &"� `��M9��7�Q�NzJ�?�@}TUb�7R����{62Z ��>�ҵ�d��;���
9��M<��0���N^ڏO�2�'����'(�/��@VR��nժs{�����3nU)�L1/O�DQQ�h��r��0�D��Ѫ�o����|�ꮅ���T�Gc�S>G��{1R����
�Q�K`���6o�� �l]����V����\x�����8��;�+bR��=�\�~8ϤO_�Vcm�����D*��NI��� �)I������]D���>�$˙w����NG�C�8���%��Ϛ`]����o�p}��3}<s䘧Ȋ3��51W��@�$����&�a��]��R��`����8�f��6��9�����ox��E>��ఘ�5Y�~(�\ݤ���σn�	y���lo,GZP�"t#Q&��P\V�[l;��,>a+a1��t� ��^��7�Mt\�5�H��`�K����%������ޝ-T��d۟������9̸�s
���lzE�X�{�#w���̡l��{� !���D9k��Ի^YUKv�B$ �Re�P{�$`�)��Qr�(&d
�rO��{ac�d���ꪮ�!
��G=�TY��IWu-��P���`=a��Q���F
�8s1!�&|$?	t�Ʉ�(�#�q'����fM��[�nқ�0��WHf�Zt���ĩ 2�xH�ˉU��?PK   �I~X=���  l     jsons/user_defined.json���n�0E%�Z$8|��]E)�>V�Q�"�P(��j���T'�.�$r��rx/�C��5h����_�T������6.lPB	��nX��Z����������[��6���7��߆2�#0o�/�U���FBe�R�Qi�He�W���Tdh��Qϱu����*X������ޔ=�2OZ��Z��\ՠ���ii��V�ۦGD 	���P����ٌ{)R;���3�N��0�����(���a���D�@!I^P9�m������'��ڌh��f�l!ΰ+Uw1p>��G:�K��|.]^�Ϟ\;;w����8���X�K�i���s�ư����ң�i2?�dFSSԬq�r�����0^g�2�Y���G�S�D���`r�%���`r2��"M��/����:$�^��v�������|��bon꿇fc|���VLS0�T���r��R�ʅ����s���0���N�(� ��}9*D�0�����G��^Ȃ�!��F�`���?PK
   �I~X;H)  h�                   cirkitFile.jsonPK
   �ZzX���7)� 
� /             V  images/0da2d01e-ca13-4f8a-b549-f8454ec0f5dd.pngPK
   2acX�#�(~ I� /             � images/e51fe3aa-205e-4659-a3a1-ad304791dd1d.pngPK
   �YzX؞�~O7  )8  /             A� images/ea12a0eb-7632-4157-afc7-05122dfed1cd.pngPK
   �I~X=���  l               ݽ jsons/user_defined.jsonPK      �  �   